CC_L1L2LL4.bsv