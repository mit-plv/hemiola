import Vector::*;
import BuildVector::*;
import FIFO::*;
import FIFOF::*;
import RWBramCore::*;
import SpecialFIFOs::*;
import HCCIfc::*;

interface CC;
    interface Vector#(L1Num, MemRqRs#(Struct1)) l1Ifc;
    interface DMA#(Bit#(13), Struct34, Vector#(4, Bit#(64))) llDma;
endinterface

typedef struct { Bit#(6) id; Bool type_; Bit#(64) addr; Vector#(4, Bit#(64)) value;  } Struct1 deriving(Eq, Bits);
typedef struct { Bool mesi_owned; Bit#(3) mesi_status; Bit#(3) mesi_dir_st; Bit#(4) mesi_dir_sharers;  } Struct10 deriving(Eq, Bits);
typedef struct { Bit#(64) mv_addr; Struct10 mv_info;  } Struct11 deriving(Eq, Bits);
typedef struct { Struct6 lr_ir_pp; Struct9 lr_ir; Vector#(4, Bit#(64)) lr_value;  } Struct12 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(64) victim_addr; Struct10 victim_info; Vector#(4, Bit#(64)) victim_value; Struct14 victim_req;  } Struct13 deriving(Eq, Bits);
typedef struct { Bool valid; Bit#(4) data;  } Struct14 deriving(Eq, Bits);
typedef struct { Bit#(3) m_status; Struct14 m_next; Bool m_is_ul; Struct1 m_msg; Bit#(4) m_qidx; Bool m_rsb; Bit#(4) m_dl_rss_from; Bit#(4) m_dl_rss_recv; Vector#(4, Struct1) m_dl_rss;  } Struct15 deriving(Eq, Bits);
typedef struct { Bit#(3) dir_st; Bit#(2) dir_excl; Bit#(4) dir_sharers;  } Struct16 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_write; Bool info_hit; Bit#(4) info_way; Bool edir_hit; Bit#(3) edir_way; Struct5 edir_slot; Struct10 info; Bool value_write; Vector#(4, Bit#(64)) value; Struct11 may_victim; Vector#(16, Bit#(8)) reps;  } Struct17 deriving(Eq, Bits);
typedef struct { Bit#(3) victim_idx; Struct10 victim_info; Vector#(4, Bit#(64)) victim_value;  } Struct18 deriving(Eq, Bits);
typedef struct { Bit#(2) enq_type; Bit#(2) enq_ch_idx; Struct1 enq_msg;  } Struct19 deriving(Eq, Bits);
typedef struct { Struct1 in_msg; Bit#(4) in_msg_from;  } Struct2 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bool r_ul_rsb; Bit#(2) r_ul_rsbTo;  } Struct20 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bit#(4) r_dl_rss_from; Bool r_dl_rsb; Bit#(4) r_dl_rsbTo;  } Struct21 deriving(Eq, Bits);
typedef struct { Bit#(4) cs_inds; Struct1 cs_msg;  } Struct22 deriving(Eq, Bits);
typedef struct { Bit#(4) cidx; Struct1 msg;  } Struct23 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bit#(4) r_dl_rss_from;  } Struct24 deriving(Eq, Bits);
typedef struct { Bit#(64) victim_addr; Bit#(4) victim_req;  } Struct25 deriving(Eq, Bits);
typedef struct { Bit#(50) tag; Struct10 value;  } Struct26 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(4) tm_way; Struct10 tm_value;  } Struct27 deriving(Eq, Bits);
typedef struct { Bit#(50) tag; Struct29 value;  } Struct28 deriving(Eq, Bits);
typedef struct { Bool mesi_edir_owned; Bit#(3) mesi_edir_st; Bit#(4) mesi_edir_sharers;  } Struct29 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Struct1 r_msg; Bit#(4) r_msg_from;  } Struct3 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(3) tm_way; Struct29 tm_value;  } Struct30 deriving(Eq, Bits);
typedef struct { Bit#(9) addr; Struct26 datain;  } Struct31 deriving(Eq, Bits);
typedef struct { Bit#(1) acc_type; Vector#(16, Bit#(8)) acc_reps; Bit#(9) acc_index; Bit#(4) acc_way;  } Struct32 deriving(Eq, Bits);
typedef struct { Bit#(9) addr; Struct28 datain;  } Struct33 deriving(Eq, Bits);
typedef struct { Bit#(13) addr; Vector#(4, Bit#(64)) datain;  } Struct34 deriving(Eq, Bits);
typedef struct { Bool valid; Struct13 data;  } Struct35 deriving(Eq, Bits);
typedef struct { Bit#(9) addr; Vector#(16, Bit#(8)) datain;  } Struct36 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Struct1 r_msg; Bit#(4) r_msg_from;  } Struct37 deriving(Eq, Bits);
typedef struct { Bool s_has_slot; Bool s_conflict; Bit#(3) s_id;  } Struct38 deriving(Eq, Bits);
typedef struct { Bool valid; Bit#(2) data;  } Struct39 deriving(Eq, Bits);
typedef struct { Bool s_has_slot; Bool s_conflict; Bit#(4) s_id;  } Struct4 deriving(Eq, Bits);
typedef struct { Bool ir_is_rs_rel; Struct1 ir_msg; Bit#(4) ir_msg_from; Bit#(3) ir_mshr_id; Struct39 ir_by_victim;  } Struct40 deriving(Eq, Bits);
typedef struct { Bit#(8) info_index; Bool info_hit; Bit#(2) info_way; Bool edir_hit; void edir_way; Struct42 edir_slot; Struct10 info; Struct11 may_victim; Vector#(4, Bit#(8)) reps;  } Struct41 deriving(Eq, Bits);
typedef struct { Bool valid; void data;  } Struct42 deriving(Eq, Bits);
typedef struct { Struct40 lr_ir_pp; Struct41 lr_ir; Vector#(4, Bit#(64)) lr_value;  } Struct43 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(64) victim_addr; Struct10 victim_info; Vector#(4, Bit#(64)) victim_value; Struct5 victim_req;  } Struct44 deriving(Eq, Bits);
typedef struct { Bit#(3) m_status; Struct5 m_next; Bool m_is_ul; Struct1 m_msg; Bit#(4) m_qidx; Bool m_rsb; Bit#(4) m_dl_rss_from; Bit#(4) m_dl_rss_recv; Vector#(4, Struct1) m_dl_rss;  } Struct45 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_write; Bool info_hit; Bit#(2) info_way; Bool edir_hit; void edir_way; Struct42 edir_slot; Struct10 info; Bool value_write; Vector#(4, Bit#(64)) value; Struct11 may_victim; Vector#(4, Bit#(8)) reps;  } Struct46 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bool r_ul_rsb; Bit#(2) r_ul_rsbTo;  } Struct47 deriving(Eq, Bits);
typedef struct { Bit#(2) victim_idx; Struct10 victim_info; Vector#(4, Bit#(64)) victim_value;  } Struct48 deriving(Eq, Bits);
typedef struct { Bit#(64) victim_addr; Bit#(3) victim_req;  } Struct49 deriving(Eq, Bits);
typedef struct { Bool valid; Bit#(3) data;  } Struct5 deriving(Eq, Bits);
typedef struct { Bit#(51) tag; Struct10 value;  } Struct50 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(2) tm_way; Struct10 tm_value;  } Struct51 deriving(Eq, Bits);
typedef struct { Bit#(8) addr; Struct50 datain;  } Struct52 deriving(Eq, Bits);
typedef struct { Bit#(1) acc_type; Vector#(4, Bit#(8)) acc_reps; Bit#(8) acc_index; Bit#(2) acc_way;  } Struct53 deriving(Eq, Bits);
typedef struct { Bit#(10) addr; Vector#(4, Bit#(64)) datain;  } Struct54 deriving(Eq, Bits);
typedef struct { Bool valid; Struct44 data;  } Struct55 deriving(Eq, Bits);
typedef struct { Bit#(8) addr; Vector#(4, Bit#(8)) datain;  } Struct56 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bit#(4) r_dl_rss_from; Bool r_dl_rsb; Bit#(4) r_dl_rsbTo;  } Struct57 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bit#(4) r_dl_rss_from;  } Struct58 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bit#(64) r_addr;  } Struct59 deriving(Eq, Bits);
typedef struct { Bool ir_is_rs_rel; Struct1 ir_msg; Bit#(4) ir_msg_from; Bit#(4) ir_mshr_id; Struct5 ir_by_victim;  } Struct6 deriving(Eq, Bits);
typedef struct { Bit#(2) r_midx; Struct1 r_msg;  } Struct7 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bit#(64) r_addr;  } Struct8 deriving(Eq, Bits);
typedef struct { Bit#(9) info_index; Bool info_hit; Bit#(4) info_way; Bool edir_hit; Bit#(3) edir_way; Struct5 edir_slot; Struct10 info; Struct11 may_victim; Vector#(16, Bit#(8)) reps;  } Struct9 deriving(Eq, Bits);

interface Module1;
    method Action enq_fifoCRqInput_00 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput_00 ();
endinterface

module mkModule1
    (Module1);
    Reg#(Vector#(4, Struct2)) elt_fifoCRqInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoCRqInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoCRqInput_00 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoCRqInput_00 <- mkReg(True);
    Reg#(Bool) full_fifoCRqInput_00 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoCRqInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoCRqInput_00 <- mkReg(unpack(0));

    rule count_fifoCRqInput_00;

        let x_0 = (countDone_fifoCRqInput_00);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoCRqInput_00);
        counter_fifoCRqInput_00 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoCRqInput_00);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoCRqInput_00);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoCRqInput_00:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoCRqInput_00:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoCRqInput_00:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoCRqInput_00:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoCRqInput_00 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoCRqInput_00 (Struct2 x_0);
        let x_1 = (full_fifoCRqInput_00);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_00);
        let x_3 = (enqP_fifoCRqInput_00);
        let x_4 = (deqP_fifoCRqInput_00);
        elt_fifoCRqInput_00 <= update (x_2, x_3, x_0);
        empty_fifoCRqInput_00 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoCRqInput_00 <= (x_4) == (x_5);
        enqP_fifoCRqInput_00 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput_00 ();
        let x_1 = (empty_fifoCRqInput_00);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_00);
        let x_3 = (enqP_fifoCRqInput_00);
        let x_4 = (deqP_fifoCRqInput_00);
        full_fifoCRqInput_00 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoCRqInput_00 <= (x_3) == (x_5);
        deqP_fifoCRqInput_00 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module2;
    method Action enq_fifoCRsInput_00 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRsInput_00 ();
endinterface

module mkModule2
    (Module2);
    Reg#(Vector#(4, Struct2)) elt_fifoCRsInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoCRsInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoCRsInput_00 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoCRsInput_00 <- mkReg(True);
    Reg#(Bool) full_fifoCRsInput_00 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoCRsInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoCRsInput_00 <- mkReg(unpack(0));

    rule count_fifoCRsInput_00;

        let x_0 = (countDone_fifoCRsInput_00);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoCRsInput_00);
        counter_fifoCRsInput_00 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoCRsInput_00);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoCRsInput_00);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoCRsInput_00:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoCRsInput_00:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoCRsInput_00:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoCRsInput_00:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoCRsInput_00 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoCRsInput_00 (Struct2 x_0);
        let x_1 = (full_fifoCRsInput_00);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRsInput_00);
        let x_3 = (enqP_fifoCRsInput_00);
        let x_4 = (deqP_fifoCRsInput_00);
        elt_fifoCRsInput_00 <= update (x_2, x_3, x_0);
        empty_fifoCRsInput_00 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoCRsInput_00 <= (x_4) == (x_5);
        enqP_fifoCRsInput_00 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoCRsInput_00 ();
        let x_1 = (empty_fifoCRsInput_00);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRsInput_00);
        let x_3 = (enqP_fifoCRsInput_00);
        let x_4 = (deqP_fifoCRsInput_00);
        full_fifoCRsInput_00 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoCRsInput_00 <= (x_3) == (x_5);
        deqP_fifoCRsInput_00 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module3;
    method Action enq_fifoPInput_00 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoPInput_00 ();
endinterface

module mkModule3
    (Module3);
    Reg#(Vector#(4, Struct2)) elt_fifoPInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoPInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoPInput_00 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoPInput_00 <- mkReg(True);
    Reg#(Bool) full_fifoPInput_00 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoPInput_00 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoPInput_00 <- mkReg(unpack(0));

    rule count_fifoPInput_00;

        let x_0 = (countDone_fifoPInput_00);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoPInput_00);
        counter_fifoPInput_00 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoPInput_00);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoPInput_00);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoPInput_00:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoPInput_00:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoPInput_00:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoPInput_00:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoPInput_00 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoPInput_00 (Struct2 x_0);
        let x_1 = (full_fifoPInput_00);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_00);
        let x_3 = (enqP_fifoPInput_00);
        let x_4 = (deqP_fifoPInput_00);
        elt_fifoPInput_00 <= update (x_2, x_3, x_0);
        empty_fifoPInput_00 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoPInput_00 <= (x_4) == (x_5);
        enqP_fifoPInput_00 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoPInput_00 ();
        let x_1 = (empty_fifoPInput_00);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_00);
        let x_3 = (enqP_fifoPInput_00);
        let x_4 = (deqP_fifoPInput_00);
        full_fifoPInput_00 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoPInput_00 <= (x_3) == (x_5);
        deqP_fifoPInput_00 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module4;
    method Action enq_fifoN2I_00 (Struct6 x_0);
    method ActionValue#(Struct6) deq_fifoN2I_00 ();
endinterface

module mkModule4
    (Module4);
    Reg#(Struct6) elt_fifoN2I_00 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoN2I_00 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoN2I_00 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoN2I_00 <- mkReg(unpack(0));

    rule count_fifoN2I_00;

        let x_0 = (countDone_fifoN2I_00);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoN2I_00);
        counter_fifoN2I_00 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoN2I_00);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoN2I_00);
            $display ("-- IR fifoN2I_00: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoN2I_00 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoN2I_00 (Struct6 x_0);
        let x_1 = (full_fifoN2I_00);
        when (! (x_1), noAction);
        elt_fifoN2I_00 <= x_0;
        full_fifoN2I_00 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct6) deq_fifoN2I_00 ();
        let x_1 = (full_fifoN2I_00);
        when (x_1, noAction);
        let x_2 = (elt_fifoN2I_00);
        full_fifoN2I_00 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module5;
    method Action enq_fifoI2L_00 (Struct6 x_0);
    method ActionValue#(Struct6) deq_fifoI2L_00 ();
endinterface

module mkModule5
    (Module5);
    Reg#(Struct6) elt_fifoI2L_00 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoI2L_00 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoI2L_00 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoI2L_00 <- mkReg(unpack(0));

    rule count_fifoI2L_00;

        let x_0 = (countDone_fifoI2L_00);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoI2L_00);
        counter_fifoI2L_00 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoI2L_00);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoI2L_00);
            $display ("-- IR fifoI2L_00: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoI2L_00 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoI2L_00 (Struct6 x_0);
        let x_1 = (full_fifoI2L_00);
        when (! (x_1), noAction);
        elt_fifoI2L_00 <= x_0;
        full_fifoI2L_00 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct6) deq_fifoI2L_00 ();
        let x_1 = (full_fifoI2L_00);
        when (x_1, noAction);
        let x_2 = (elt_fifoI2L_00);
        full_fifoI2L_00 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module6;
    method Action enq_fifoL2E_00 (Struct12 x_0);
    method ActionValue#(Struct12) deq_fifoL2E_00 ();
endinterface

module mkModule6
    (Module6);
    Reg#(Struct12) elt_fifoL2E_00 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoL2E_00 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoL2E_00 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoL2E_00 <- mkReg(unpack(0));

    rule count_fifoL2E_00;

        let x_0 = (countDone_fifoL2E_00);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoL2E_00);
        counter_fifoL2E_00 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoL2E_00);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoL2E_00);
            $display ("-- LR fifoL2E_00: %b %x %b %x %x %x %b %x %x %b %x %b %x %b %x", ((x_3).lr_ir_pp).ir_is_rs_rel, (((x_3).lr_ir_pp).ir_msg).id, (((x_3).lr_ir_pp).ir_msg).type_, (((x_3).lr_ir_pp).ir_msg).addr, ((x_3).lr_ir_pp).ir_msg_from, ((x_3).lr_ir_pp).ir_mshr_id, (((x_3).lr_ir_pp).ir_by_victim).valid, (((x_3).lr_ir_pp).ir_by_victim).data, ((x_3).lr_ir).info_index, ((x_3).lr_ir).info_hit, ((x_3).lr_ir).info_way, ((x_3).lr_ir).edir_hit, ((x_3).lr_ir).edir_way, (((x_3).lr_ir).edir_slot).valid, (((x_3).lr_ir).edir_slot).data);
            countDone_fifoL2E_00 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoL2E_00 (Struct12 x_0);
        let x_1 = (full_fifoL2E_00);
        when (! (x_1), noAction);
        elt_fifoL2E_00 <= x_0;
        full_fifoL2E_00 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct12) deq_fifoL2E_00 ();
        let x_1 = (full_fifoL2E_00);
        when (x_1, noAction);
        let x_2 = (elt_fifoL2E_00);
        full_fifoL2E_00 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module7;
    method ActionValue#(Struct5) victims__00__findVictim (Bit#(64) x_0);
    method ActionValue#(Struct13) victims__00__getVictim (Bit#(3) x_0);
    method Action victims__00__setVictim (Struct18 x_0);
    method Action victims__00__registerVictim (Struct13 x_0);
    method ActionValue#(Struct13) victims__00__getFirstVictim ();
    method ActionValue#(Bool) victims__00__hasVictim ();
    method Action victims__00__setVictimRq (Struct25 x_0);
    method ActionValue#(Bit#(4)) victims__00__releaseVictim (Bit#(64) x_0);
endinterface

module mkModule7
    (Module7);
    Reg#(Vector#(8, Struct13)) victimRegs__00 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct5) victims__00__findVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__00);
        Struct13 x_2 =
        ((x_1)[(Bit#(3))'(3'h0)]);
        let x_17 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            x_17 = Struct5 {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)};
        end else begin
            Struct13 x_3 =
            ((x_1)[(Bit#(3))'(3'h1)]);
            let x_16 = ?;
            if (((x_3).victim_valid) && (((x_3).victim_addr) == (x_0)))
                begin
                x_16 = Struct5 {valid : (Bool)'(True), data :
                (Bit#(3))'(3'h1)};
            end else begin
                Struct13 x_4 =
                ((x_1)[(Bit#(3))'(3'h2)]);
                let x_15 = ?;
                if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                    begin
                    x_15 = Struct5 {valid : (Bool)'(True), data :
                    (Bit#(3))'(3'h2)};
                end else begin
                    Struct13 x_5 =
                    ((x_1)[(Bit#(3))'(3'h3)]);
                    let x_14 = ?;
                    if (((x_5).victim_valid) && (((x_5).victim_addr) ==
                        (x_0))) begin
                        x_14 = Struct5 {valid : (Bool)'(True), data :
                        (Bit#(3))'(3'h3)};
                    end else begin
                        Struct13 x_6 =
                        ((x_1)[(Bit#(3))'(3'h4)]);
                        let x_13 = ?;
                        if (((x_6).victim_valid) && (((x_6).victim_addr) ==
                            (x_0))) begin
                            x_13 = Struct5 {valid : (Bool)'(True), data :
                            (Bit#(3))'(3'h4)};
                        end else begin
                            Struct13 x_7 =
                            ((x_1)[(Bit#(3))'(3'h5)]);
                            let x_12 = ?;
                            if (((x_7).victim_valid) && (((x_7).victim_addr)
                                == (x_0))) begin
                                x_12 = Struct5 {valid : (Bool)'(True), data :
                                (Bit#(3))'(3'h5)};
                            end else begin
                                Struct13 x_8 =
                                ((x_1)[(Bit#(3))'(3'h6)]);
                                let x_11 = ?;
                                if (((x_8).victim_valid) &&
                                    (((x_8).victim_addr) == (x_0))) begin
                                    x_11 = Struct5 {valid : (Bool)'(True),
                                    data : (Bit#(3))'(3'h6)};
                                end else begin
                                    Struct13 x_9 =
                                    ((x_1)[(Bit#(3))'(3'h7)]);
                                    let x_10 = ?;
                                    if (((x_9).victim_valid) &&
                                        (((x_9).victim_addr) == (x_0)))
                                        begin
                                        x_10 = Struct5 {valid :
                                        (Bool)'(True), data :
                                        (Bit#(3))'(3'h7)};
                                    end else begin
                                        x_10 = Struct5 {valid :
                                        (Bool)'(False), data : unpack(0)};
                                    end
                                    x_11 = x_10;
                                end
                                x_12 = x_11;
                            end
                            x_13 = x_12;
                        end
                        x_14 = x_13;
                    end
                    x_15 = x_14;
                end
                x_16 = x_15;
            end
            x_17 = x_16;
        end
        return x_17;
    endmethod

    method ActionValue#(Struct13) victims__00__getVictim (Bit#(3) x_0);
        let x_1 = (victimRegs__00);
        return (x_1)[x_0];
    endmethod

    method Action victims__00__setVictim (Struct18 x_0);
        let x_1 = (victimRegs__00);
        Struct13 x_2 = ((x_1)[(x_0).victim_idx]);
        Struct13 x_3 = (Struct13 {victim_valid : (Bool)'(True), victim_addr :
        (x_2).victim_addr, victim_info : (x_0).victim_info, victim_value :
        (x_0).victim_value, victim_req : (x_2).victim_req});
        victimRegs__00 <= update (x_1, (x_0).victim_idx, x_3);
    endmethod

    method Action victims__00__registerVictim (Struct13 x_0);
        let x_1 = (victimRegs__00);
        Struct5 x_2 = ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid ?
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid ?
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid ?
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid ?
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid ?
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid ?
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid ?
        ((((x_1)[(Bit#(3))'(3'h0)]).victim_valid ? (Struct5 {valid :
        (Bool)'(False), data : unpack(0)}) : (Struct5 {valid : (Bool)'(True),
        data : (Bit#(3))'(3'h0)}))) : (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}))) : (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}))) : (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}))) : (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}))) : (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}))) : (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h6)}))) : (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h7)})));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        victimRegs__00 <= update (x_1, x_3, x_0);
    endmethod

    method ActionValue#(Struct13) victims__00__getFirstVictim ();
        let x_1 = (victimRegs__00);
        Struct35 x_2 = (((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h7)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h7)]}) :
        (((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h6)]}) :
        (((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h5)]}) :
        (((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h4)]}) :
        (((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h3)]}) :
        (((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h2)]}) :
        (((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h1)]}) :
        (((((x_1)[(Bit#(3))'(3'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).victim_req).valid)) ? (Struct35 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h0)]}) : (Struct35 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method ActionValue#(Bool) victims__00__hasVictim ();
        let x_1 = (victimRegs__00);
        Bool x_2 = (((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h7)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(3))'(3'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).victim_req).valid)) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))))))))))));
        return x_2;
    endmethod

    method Action victims__00__setVictimRq (Struct25 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(4) x_2 = ((x_0).victim_req);
        let x_3 = (victimRegs__00);
        Struct13 x_4 =
        ((x_3)[(Bit#(3))'(3'h7)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct13 x_5 = (Struct13 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct14 {valid :
            (Bool)'(True), data : x_2}});
            victimRegs__00 <= update (x_3, (Bit#(3))'(3'h7), x_5);
        end else begin
            Struct13 x_6 =
            ((x_3)[(Bit#(3))'(3'h6)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct13 x_7 = (Struct13 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct14 {valid : (Bool)'(True), data :
                x_2}});
                victimRegs__00 <= update (x_3, (Bit#(3))'(3'h6), x_7);
            end else begin
                Struct13 x_8 =
                ((x_3)[(Bit#(3))'(3'h5)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct13 x_9 = (Struct13 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct14 {valid :
                    (Bool)'(True), data : x_2}});
                    victimRegs__00 <= update (x_3, (Bit#(3))'(3'h5), x_9);
                end else begin
                    Struct13 x_10 =
                    ((x_3)[(Bit#(3))'(3'h4)]);
                    if (((x_10).victim_valid) && (((x_10).victim_addr) ==
                        (x_1))) begin
                        Struct13 x_11 = (Struct13 {victim_valid :
                        (x_10).victim_valid, victim_addr :
                        (x_10).victim_addr, victim_info : (x_10).victim_info,
                        victim_value : (x_10).victim_value, victim_req :
                        Struct14 {valid : (Bool)'(True), data :
                        x_2}});
                        victimRegs__00 <= update (x_3, (Bit#(3))'(3'h4),
                        x_11);
                    end else begin
                        Struct13 x_12 =
                        ((x_3)[(Bit#(3))'(3'h3)]);
                        if (((x_12).victim_valid) && (((x_12).victim_addr) ==
                            (x_1))) begin
                            Struct13 x_13 = (Struct13 {victim_valid :
                            (x_12).victim_valid, victim_addr :
                            (x_12).victim_addr, victim_info :
                            (x_12).victim_info, victim_value :
                            (x_12).victim_value, victim_req : Struct14 {valid
                            : (Bool)'(True), data : x_2}});
                            victimRegs__00 <= update (x_3, (Bit#(3))'(3'h3),
                            x_13);
                        end else begin
                            Struct13 x_14 =
                            ((x_3)[(Bit#(3))'(3'h2)]);
                            if (((x_14).victim_valid) &&
                                (((x_14).victim_addr) == (x_1)))
                                begin
                                Struct13 x_15 = (Struct13 {victim_valid :
                                (x_14).victim_valid, victim_addr :
                                (x_14).victim_addr, victim_info :
                                (x_14).victim_info, victim_value :
                                (x_14).victim_value, victim_req : Struct14
                                {valid : (Bool)'(True), data :
                                x_2}});
                                victimRegs__00 <= update (x_3,
                                (Bit#(3))'(3'h2), x_15);
                            end else begin
                                Struct13 x_16 =
                                ((x_3)[(Bit#(3))'(3'h1)]);
                                if (((x_16).victim_valid) &&
                                    (((x_16).victim_addr) == (x_1)))
                                    begin
                                    Struct13 x_17 = (Struct13 {victim_valid :
                                    (x_16).victim_valid, victim_addr :
                                    (x_16).victim_addr, victim_info :
                                    (x_16).victim_info, victim_value :
                                    (x_16).victim_value, victim_req :
                                    Struct14 {valid : (Bool)'(True), data :
                                    x_2}});
                                    victimRegs__00 <= update (x_3,
                                    (Bit#(3))'(3'h1), x_17);
                                end else begin
                                    Struct13 x_18 =
                                    ((x_3)[(Bit#(3))'(3'h0)]);
                                    if (((x_18).victim_valid) &&
                                        (((x_18).victim_addr) == (x_1)))
                                        begin
                                        Struct13 x_19 = (Struct13
                                        {victim_valid : (x_18).victim_valid,
                                        victim_addr : (x_18).victim_addr,
                                        victim_info : (x_18).victim_info,
                                        victim_value : (x_18).victim_value,
                                        victim_req : Struct14 {valid :
                                        (Bool)'(True), data :
                                        x_2}});
                                        victimRegs__00 <= update (x_3,
                                        (Bit#(3))'(3'h0), x_19);
                                    end else begin

                                    end
                                end
                            end
                        end
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Bit#(4)) victims__00__releaseVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__00);
        Struct13 x_2 =
        ((x_1)[(Bit#(3))'(3'h0)]);
        let x_25 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victimRegs__00 <= update (x_1, (Bit#(3))'(3'h0),
            unpack(0));
            Bit#(4) x_3 = (((x_2).victim_req).data);
            x_25 = x_3;
        end else begin
            Struct13 x_4 =
            ((x_1)[(Bit#(3))'(3'h1)]);
            let x_24 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victimRegs__00 <= update (x_1, (Bit#(3))'(3'h1),
                unpack(0));
                Bit#(4) x_5 = (((x_4).victim_req).data);
                x_24 = x_5;
            end else begin
                Struct13 x_6 =
                ((x_1)[(Bit#(3))'(3'h2)]);
                let x_23 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victimRegs__00 <= update (x_1, (Bit#(3))'(3'h2),
                    unpack(0));
                    Bit#(4) x_7 = (((x_6).victim_req).data);
                    x_23 = x_7;
                end else begin
                    Struct13 x_8 =
                    ((x_1)[(Bit#(3))'(3'h3)]);
                    let x_22 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victimRegs__00 <= update (x_1, (Bit#(3))'(3'h3),
                        unpack(0));
                        Bit#(4) x_9 = (((x_8).victim_req).data);
                        x_22 = x_9;
                    end else begin
                        Struct13 x_10 =
                        ((x_1)[(Bit#(3))'(3'h4)]);
                        let x_21 = ?;
                        if (((x_10).victim_valid) && (((x_10).victim_addr) ==
                            (x_0))) begin
                            victimRegs__00 <= update (x_1, (Bit#(3))'(3'h4),
                            unpack(0));
                            Bit#(4) x_11 = (((x_10).victim_req).data);
                            x_21 = x_11;
                        end else begin
                            Struct13 x_12 =
                            ((x_1)[(Bit#(3))'(3'h5)]);
                            let x_20 = ?;
                            if (((x_12).victim_valid) &&
                                (((x_12).victim_addr) == (x_0)))
                                begin
                                victimRegs__00 <= update (x_1,
                                (Bit#(3))'(3'h5), unpack(0));
                                Bit#(4) x_13 =
                                (((x_12).victim_req).data);
                                x_20 = x_13;
                            end else begin
                                Struct13 x_14 =
                                ((x_1)[(Bit#(3))'(3'h6)]);
                                let x_19 = ?;
                                if (((x_14).victim_valid) &&
                                    (((x_14).victim_addr) == (x_0)))
                                    begin
                                    victimRegs__00 <= update (x_1,
                                    (Bit#(3))'(3'h6), unpack(0));
                                    Bit#(4) x_15 =
                                    (((x_14).victim_req).data);
                                    x_19 = x_15;
                                end else begin
                                    Struct13 x_16 =
                                    ((x_1)[(Bit#(3))'(3'h7)]);
                                    let x_18 = ?;
                                    if (((x_16).victim_valid) &&
                                        (((x_16).victim_addr) == (x_0)))
                                        begin
                                        victimRegs__00 <= update (x_1,
                                        (Bit#(3))'(3'h7), unpack(0));
                                        Bit#(4) x_17 =
                                        (((x_16).victim_req).data);
                                        x_18 = x_17;
                                    end else begin
                                        x_18 = unpack(0);
                                    end
                                    x_19 = x_18;
                                end
                                x_20 = x_19;
                            end
                            x_21 = x_20;
                        end
                        x_22 = x_21;
                    end
                    x_23 = x_22;
                end
                x_24 = x_23;
            end
            x_25 = x_24;
        end
        return x_25;
    endmethod
endmodule

interface Module8;
    method Action rdReq_infoRam__00__15 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__15 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__15 ();
endinterface

module mkModule8 (Module8);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h1f, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__15 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__15 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__15 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module9;
    method Action rdReq_infoRam__00__14 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__14 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__14 ();
endinterface

module mkModule9 (Module9);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h1e, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__14 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__14 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__14 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module10;
    method Action rdReq_infoRam__00__13 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__13 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__13 ();
endinterface

module mkModule10 (Module10);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h1d, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__13 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__13 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__13 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module11;
    method Action rdReq_infoRam__00__12 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__12 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__12 ();
endinterface

module mkModule11 (Module11);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h1c, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__12 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__12 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__12 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module12;
    method Action rdReq_infoRam__00__11 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__11 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__11 ();
endinterface

module mkModule12 (Module12);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h1b, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__11 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__11 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__11 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module13;
    method Action rdReq_infoRam__00__10 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__10 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__10 ();
endinterface

module mkModule13 (Module13);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h1a, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__10 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__10 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__10 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module14;
    method Action rdReq_infoRam__00__9 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__9 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__9 ();
endinterface

module mkModule14 (Module14);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h19, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__9 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__9 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__9 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module15;
    method Action rdReq_infoRam__00__8 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__8 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__8 ();
endinterface

module mkModule15 (Module15);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h18, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__8 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__8 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__8 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module16;
    method Action rdReq_infoRam__00__7 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__7 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__7 ();
endinterface

module mkModule16 (Module16);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h17, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__7 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__7 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__7 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module17;
    method Action rdReq_infoRam__00__6 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__6 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__6 ();
endinterface

module mkModule17 (Module17);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h16, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__6 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__6 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__6 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module18;
    method Action rdReq_infoRam__00__5 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__5 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__5 ();
endinterface

module mkModule18 (Module18);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h15, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__5 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__5 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__5 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module19;
    method Action rdReq_infoRam__00__4 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__4 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__4 ();
endinterface

module mkModule19 (Module19);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h14, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__4 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__4 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__4 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module20;
    method Action rdReq_infoRam__00__3 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__3 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__3 ();
endinterface

module mkModule20 (Module20);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h13, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__3 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__3 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module21;
    method Action rdReq_infoRam__00__2 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__2 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__2 ();
endinterface

module mkModule21 (Module21);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h12, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__2 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__2 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module22;
    method Action rdReq_infoRam__00__1 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__1 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__1 ();
endinterface

module mkModule22 (Module22);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h11, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__1 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__1 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module23;
    method Action rdReq_infoRam__00__0 (Bit#(9) x_0);
    method Action wrReq_infoRam__00__0 (Struct31 x_0);
    method ActionValue#(Struct26) rdResp_infoRam__00__0 ();
endinterface

module mkModule23 (Module23);
    RWBramCore#(Bit#(9), Struct26) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct26 {tag: 50'h10, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__0 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__0 (Struct31 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct26) rdResp_infoRam__00__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module24;
    method Action rdReq_edirRam__00__7 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__7 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__7 ();
endinterface

module mkModule24 (Module24);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h27, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__7 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__7 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__7 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module25;
    method Action rdReq_edirRam__00__6 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__6 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__6 ();
endinterface

module mkModule25 (Module25);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h26, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__6 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__6 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__6 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module26;
    method Action rdReq_edirRam__00__5 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__5 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__5 ();
endinterface

module mkModule26 (Module26);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h25, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__5 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__5 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__5 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module27;
    method Action rdReq_edirRam__00__4 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__4 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__4 ();
endinterface

module mkModule27 (Module27);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h24, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__4 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__4 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__4 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module28;
    method Action rdReq_edirRam__00__3 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__3 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__3 ();
endinterface

module mkModule28 (Module28);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h23, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__3 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__3 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module29;
    method Action rdReq_edirRam__00__2 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__2 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__2 ();
endinterface

module mkModule29 (Module29);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h22, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__2 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__2 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module30;
    method Action rdReq_edirRam__00__1 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__1 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__1 ();
endinterface

module mkModule30 (Module30);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h21, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__1 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__1 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module31;
    method Action rdReq_edirRam__00__0 (Bit#(9) x_0);
    method Action wrReq_edirRam__00__0 (Struct33 x_0);
    method ActionValue#(Struct28) rdResp_edirRam__00__0 ();
endinterface

module mkModule31 (Module31);
    RWBramCore#(Bit#(9), Struct28) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct28 {tag: 50'h20, value: Struct29 {mesi_edir_owned: False, mesi_edir_st: 3'h1, mesi_edir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__0 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__0 (Struct33 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct28) rdResp_edirRam__00__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module32;
    method Action rdReq_dataRam__00 (Bit#(13) x_0);
    method Action wrReq_dataRam__00 (Struct34 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__00 ();
endinterface

module mkModule32 (Module32);
    RWBramCore#(Bit#(13), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(13)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__00 (Bit#(13) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__00 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__00 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module33;
    method Action rdReq_repRam__00 (Bit#(9) x_0);
    method Action wrReq_repRam__00 (Struct36 x_0);
    method ActionValue#(Vector#(16, Bit#(8))) rdResp_repRam__00 ();
endinterface

module mkModule33 (Module33);
    RWBramCore#(Bit#(9), Vector#(16, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1, 8'h1);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__00 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__00 (Struct36 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(16, Bit#(8))) rdResp_repRam__00 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module34;
    method ActionValue#(Struct15) getMSHR_00 (Bit#(4) x_0);
    method ActionValue#(Struct4) getPRqSlot_00 (Struct3 x_0);
    method ActionValue#(Struct4) getCRqSlot_00 (Struct3 x_0);
    method ActionValue#(Struct3) getWait_00 ();
    method Action registerUL_00 (Struct20 x_0);
    method Action registerDL_00 (Struct21 x_0);
    method Action canImm_00 (Bit#(64) x_0);
    method ActionValue#(Bit#(4)) setULImm_00 (Struct1 x_0);
    method Action transferUpDown_00 (Struct24 x_0);
    method Action addRs_00 (Struct7 x_0);
    method ActionValue#(Bit#(4)) getULReady_00 (Bit#(64) x_0);
    method ActionValue#(Struct8) getDLReady_00 ();
    method Action startRelease_00 (Bit#(4) x_0);
    method Action releaseMSHR_00 (Bit#(4) x_0);
endinterface

module mkModule34
    (Module34);
    Reg#(Vector#(12, Struct15)) rqs_00 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct15) getMSHR_00 (Bit#(4) x_0);
        let x_1 = (rqs_00);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct4) getPRqSlot_00 (Struct3 x_0);
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        || (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : ((Bool)'(False))))))))))))))))))))))))));
        Struct14 x_7 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) :
        (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) :
        (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) :
        (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) :
        (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) :
        (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        Bool x_8 = ((x_7).valid);
        Struct4 x_9 = (Struct4 {s_has_slot : (x_3) && (! (x_6)), s_conflict :
        x_8, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(12, Struct15) x_10 = (update (x_1, x_4, Struct15
            {m_status : (x_8 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))),
            m_next : Struct14 {valid : (Bool)'(False), data : unpack(0)},
            m_is_ul : unpack(0), m_msg : (x_0).r_msg, m_qidx :
            (x_0).r_msg_from, m_rsb : unpack(0), m_dl_rss_from : unpack(0),
            m_dl_rss_recv : unpack(0), m_dl_rss :
            unpack(0)}));
            let x_14 = ?;
            if (x_8) begin
                Bit#(4) x_11 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
                ((Bit#(3))'(3'h0)))) && (!
                ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h0)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h1)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h2)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h3)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h4)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h5)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h6)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h7)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h8)) : ((((!
                ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'h9)) : ((((!
                ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'ha)) : ((((!
                ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
                (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ?
                ((Bit#(4))'(4'hb)) :
                (unpack(0))))))))))))))))))))))))));
                Struct15 x_12 = ((x_1)[x_11]);
                Vector#(12, Struct15) x_13 = (update (x_10, x_11, Struct15
                {m_status : (x_12).m_status, m_next : (x_8 ? (Struct14 {valid
                : (Bool)'(True), data : x_4}) : ((x_12).m_next)), m_is_ul :
                (x_12).m_is_ul, m_msg : (x_12).m_msg, m_qidx : (x_12).m_qidx,
                m_rsb : (x_12).m_rsb, m_dl_rss_from : (x_12).m_dl_rss_from,
                m_dl_rss_recv : (x_12).m_dl_rss_recv, m_dl_rss :
                (x_12).m_dl_rss}));
                x_14 = x_13;
            end else begin
                x_14 = x_10;
            end
            rqs_00 <= x_14;
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct4) getCRqSlot_00 (Struct3 x_0);
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))))))))))))))));
        Struct14 x_7 = (((((! ((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))));
        Struct14 x_8 = (((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : (((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        Bool x_9 = ((x_7).valid);
        Bool x_10 = ((x_8).valid);
        Bool x_11 = ((x_9) || (x_10));
        Struct4 x_12 = (Struct4 {s_has_slot : (x_3) && (! (x_6)), s_conflict
        : x_11, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(12, Struct15) x_13 = (update (x_1, x_4, Struct15
            {m_status : (x_11 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))),
            m_next : Struct14 {valid : (Bool)'(False), data : unpack(0)},
            m_is_ul : unpack(0), m_msg : (x_0).r_msg, m_qidx :
            (x_0).r_msg_from, m_rsb : unpack(0), m_dl_rss_from : unpack(0),
            m_dl_rss_recv : unpack(0), m_dl_rss :
            unpack(0)}));
            let x_17 = ?;
            if (x_11) begin
                Bit#(4) x_14 = ((x_9 ? ((x_7).data) : ((x_8).data)));
                Struct15 x_15 = ((x_1)[x_14]);
                Vector#(12, Struct15) x_16 = (update (x_13, x_14, Struct15
                {m_status : (x_15).m_status, m_next : (x_11 ? (Struct14
                {valid : (Bool)'(True), data : x_4}) : ((x_15).m_next)),
                m_is_ul : (x_15).m_is_ul, m_msg : (x_15).m_msg, m_qidx :
                (x_15).m_qidx, m_rsb : (x_15).m_rsb, m_dl_rss_from :
                (x_15).m_dl_rss_from, m_dl_rss_recv : (x_15).m_dl_rss_recv,
                m_dl_rss : (x_15).m_dl_rss}));
                x_17 = x_16;
            end else begin
                x_17 = x_13;
            end
            rqs_00 <= x_17;
        end else begin

        end
        return x_12;
    endmethod

    method ActionValue#(Struct3) getWait_00 ();
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))))))))))));
        when ((x_2).valid, noAction);
        Bit#(4) x_3 = ((x_2).data);
        Struct15 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr)[13:5]) == ((x_5)[13:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(4))'(4'h2)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr)[13:5]) == ((x_5)[13:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(4))'(4'h4)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr)[13:5]) == ((x_5)[13:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(4))'(4'h6)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr)[13:5]) == ((x_5)[13:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(4))'(4'h8)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr)[13:5]) == ((x_5)[13:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(4))'(4'ha)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr)[13:5]) == ((x_5)[13:5]))))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))))))))))))))));
        when (! (x_6), noAction);
        rqs_00 <= update (x_1, x_3, Struct15 {m_status : (Bit#(3))'(3'h4),
        m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg,
        m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : (x_4).m_dl_rss_recv, m_dl_rss :
        (x_4).m_dl_rss});
        Struct3 x_7 = (Struct3 {r_id : x_3, r_msg : (x_4).m_msg, r_msg_from :
        (x_4).m_qidx});
        return x_7;
    endmethod

    method Action registerUL_00 (Struct20 x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct15 x_3 = ((x_1)[x_2]);
        Struct15 x_4 = (Struct15 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_00 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_00 (Struct21 x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct15 x_3 = ((x_1)[x_2]);
        Struct15 x_4 = (Struct15 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_00 <= update (x_1, x_2, x_4);
    endmethod

    method Action canImm_00 (Bit#(64) x_0);
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))));
        when ((x_2).valid, noAction);
        Struct14 x_3 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        when (! ((x_3).valid), noAction);
    endmethod

    method ActionValue#(Bit#(4)) setULImm_00 (Struct1 x_0);
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))));
        when ((x_2).valid, noAction);
        Bit#(4) x_3 = ((x_2).data);
        Bit#(64) x_4 = ((x_0).addr);
        Struct14 x_5 = (((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) ==
        (x_4)) ? (Struct14 {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)})
        : (((! ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h0))))
        && (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : (((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : (((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : (((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_4)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        when (! ((x_5).valid), noAction);
        Vector#(12, Struct15) x_6 = (update (x_1, x_3, Struct15 {m_status :
        (Bit#(3))'(3'h5), m_next : Struct14 {valid : (Bool)'(False), data :
        unpack(0)}, m_is_ul : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)}));
        rqs_00 <= x_6;
        return x_3;
    endmethod

    method Action transferUpDown_00 (Struct24 x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct15 x_3 = ((x_1)[x_2]);
        Struct15 x_4 = (Struct15 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_00 <= update (x_1, x_2, x_4);
    endmethod

    method Action addRs_00 (Struct7 x_0);
        let x_1 = (rqs_00);
        Bit#(64) x_2 = (((x_0).r_msg).addr);
        Struct14 x_3 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) :
        (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) :
        (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) :
        (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) :
        (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) :
        (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_2)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        when ((x_3).valid, noAction);
        Bit#(4) x_4 = ((x_3).data);
        Struct15 x_5 = ((x_1)[x_4]);
        Struct15 x_6 = (Struct15 {m_status : (x_5).m_status, m_next :
        (x_5).m_next, m_is_ul : (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx :
        (x_5).m_qidx, m_rsb : (x_5).m_rsb, m_dl_rss_from :
        (x_5).m_dl_rss_from, m_dl_rss_recv : ((x_5).m_dl_rss_recv) |
        (((Bit#(4))'(4'h1)) << ((x_0).r_midx)), m_dl_rss : update
        ((x_5).m_dl_rss, (x_0).r_midx, (x_0).r_msg)});
        rqs_00 <= update (x_1, x_4, x_6);
    endmethod

    method ActionValue#(Bit#(4)) getULReady_00 (Bit#(64) x_0);
        let x_1 = (rqs_00);
        Bool x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)[13:5]) ==
        ((x_0)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr)[13:5]) == ((x_0)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)[13:5]) ==
        ((x_0)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr)[13:5]) == ((x_0)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)[13:5]) ==
        ((x_0)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr)[13:5]) == ((x_0)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)[13:5]) ==
        ((x_0)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr)[13:5]) == ((x_0)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)[13:5]) ==
        ((x_0)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr)[13:5]) == ((x_0)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)[13:5]) ==
        ((x_0)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr)[13:5]) == ((x_0)[13:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))))))))))))))));
        when (! (x_2), noAction);
        Struct14 x_3 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        when (! ((x_3).valid), noAction);
        Struct14 x_4 = (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) :
        (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) :
        (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) :
        (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))));
        when ((x_4).valid, noAction);
        Bit#(4) x_5 = ((x_4).data);
        return x_5;
    endmethod

    method ActionValue#(Struct8) getDLReady_00 ();
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h0)}) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h1)}) :
        (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h2)}) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h3)}) :
        (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h4)}) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h5)}) :
        (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h6)}) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h7)}) :
        (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h8)}) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'h9)}) :
        (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'ha)}) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_recv)) ? (Struct14 {valid :
        (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        when ((x_2).valid, noAction);
        Bit#(4) x_3 = ((x_2).data);
        Struct15 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr)[13:5]) ==
        ((x_5)[13:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr)[13:5]) == ((x_5)[13:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))))))))))))))));
        when (! (x_6), noAction);
        Struct8 x_7 = (Struct8 {r_id : x_3, r_addr : x_5});
        return x_7;
    endmethod

    method Action startRelease_00 (Bit#(4) x_0);
        let x_1 = (rqs_00);
        Struct15 x_2 = ((x_1)[x_0]);
        Struct15 x_3 = (Struct15 {m_status : (Bit#(3))'(3'h6), m_next :
        (x_2).m_next, m_is_ul : (x_2).m_is_ul, m_msg : (x_2).m_msg, m_qidx :
        (x_2).m_qidx, m_rsb : (x_2).m_rsb, m_dl_rss_from :
        (x_2).m_dl_rss_from, m_dl_rss_recv : (x_2).m_dl_rss_recv, m_dl_rss :
        (x_2).m_dl_rss});
        rqs_00 <= update (x_1, x_0, x_3);
    endmethod

    method Action releaseMSHR_00 (Bit#(4) x_0);
        let x_1 = (rqs_00);
        Struct15 x_2 = ((x_1)[x_0]);
        Vector#(12, Struct15) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(4) x_4 = (((x_2).m_next).data);
            Struct15 x_5 = ((x_1)[x_4]);
            Vector#(12, Struct15) x_6 = (update (x_3, x_4, Struct15 {m_status
            : (Bit#(3))'(3'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_00 <= x_7;
    endmethod
endmodule

interface Module35;
    method Action enq_fifoCRqInput_000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput_000 ();
endinterface

module mkModule35
    (Module35);
    Reg#(Vector#(4, Struct2)) elt_fifoCRqInput_000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoCRqInput_000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoCRqInput_000 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoCRqInput_000 <- mkReg(True);
    Reg#(Bool) full_fifoCRqInput_000 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoCRqInput_000 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoCRqInput_000 <- mkReg(unpack(0));

    rule count_fifoCRqInput_000;

        let x_0 = (countDone_fifoCRqInput_000);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoCRqInput_000);
        counter_fifoCRqInput_000 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoCRqInput_000);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoCRqInput_000);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoCRqInput_000:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoCRqInput_000:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoCRqInput_000:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoCRqInput_000:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoCRqInput_000 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoCRqInput_000 (Struct2 x_0);
        let x_1 = (full_fifoCRqInput_000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_000);
        let x_3 = (enqP_fifoCRqInput_000);
        let x_4 = (deqP_fifoCRqInput_000);
        elt_fifoCRqInput_000 <= update (x_2, x_3, x_0);
        empty_fifoCRqInput_000 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoCRqInput_000 <= (x_4) == (x_5);
        enqP_fifoCRqInput_000 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput_000 ();
        let x_1 = (empty_fifoCRqInput_000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_000);
        let x_3 = (enqP_fifoCRqInput_000);
        let x_4 = (deqP_fifoCRqInput_000);
        full_fifoCRqInput_000 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoCRqInput_000 <= (x_3) == (x_5);
        deqP_fifoCRqInput_000 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module36;
    method Action enq_fifoPInput_000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoPInput_000 ();
endinterface

module mkModule36
    (Module36);
    Reg#(Vector#(4, Struct2)) elt_fifoPInput_000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoPInput_000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoPInput_000 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoPInput_000 <- mkReg(True);
    Reg#(Bool) full_fifoPInput_000 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoPInput_000 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoPInput_000 <- mkReg(unpack(0));

    rule count_fifoPInput_000;

        let x_0 = (countDone_fifoPInput_000);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoPInput_000);
        counter_fifoPInput_000 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoPInput_000);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoPInput_000);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoPInput_000:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoPInput_000:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoPInput_000:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoPInput_000:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoPInput_000 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoPInput_000 (Struct2 x_0);
        let x_1 = (full_fifoPInput_000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_000);
        let x_3 = (enqP_fifoPInput_000);
        let x_4 = (deqP_fifoPInput_000);
        elt_fifoPInput_000 <= update (x_2, x_3, x_0);
        empty_fifoPInput_000 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoPInput_000 <= (x_4) == (x_5);
        enqP_fifoPInput_000 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoPInput_000 ();
        let x_1 = (empty_fifoPInput_000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_000);
        let x_3 = (enqP_fifoPInput_000);
        let x_4 = (deqP_fifoPInput_000);
        full_fifoPInput_000 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoPInput_000 <= (x_3) == (x_5);
        deqP_fifoPInput_000 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module37;
    method Action enq_fifoN2I_000 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoN2I_000 ();
endinterface

module mkModule37
    (Module37);
    Reg#(Struct40) elt_fifoN2I_000 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoN2I_000 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoN2I_000 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoN2I_000 <- mkReg(unpack(0));

    rule count_fifoN2I_000;

        let x_0 = (countDone_fifoN2I_000);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoN2I_000);
        counter_fifoN2I_000 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoN2I_000);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoN2I_000);
            $display ("-- IR fifoN2I_000: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoN2I_000 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoN2I_000 (Struct40 x_0);
        let x_1 = (full_fifoN2I_000);
        when (! (x_1), noAction);
        elt_fifoN2I_000 <= x_0;
        full_fifoN2I_000 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoN2I_000 ();
        let x_1 = (full_fifoN2I_000);
        when (x_1, noAction);
        let x_2 = (elt_fifoN2I_000);
        full_fifoN2I_000 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module38;
    method Action enq_fifoI2L_000 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoI2L_000 ();
endinterface

module mkModule38
    (Module38);
    Reg#(Struct40) elt_fifoI2L_000 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoI2L_000 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoI2L_000 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoI2L_000 <- mkReg(unpack(0));

    rule count_fifoI2L_000;

        let x_0 = (countDone_fifoI2L_000);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoI2L_000);
        counter_fifoI2L_000 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoI2L_000);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoI2L_000);
            $display ("-- IR fifoI2L_000: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoI2L_000 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoI2L_000 (Struct40 x_0);
        let x_1 = (full_fifoI2L_000);
        when (! (x_1), noAction);
        elt_fifoI2L_000 <= x_0;
        full_fifoI2L_000 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoI2L_000 ();
        let x_1 = (full_fifoI2L_000);
        when (x_1, noAction);
        let x_2 = (elt_fifoI2L_000);
        full_fifoI2L_000 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module39;
    method Action enq_fifoL2E_000 (Struct43 x_0);
    method ActionValue#(Struct43) deq_fifoL2E_000 ();
endinterface

module mkModule39
    (Module39);
    Reg#(Struct43) elt_fifoL2E_000 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoL2E_000 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoL2E_000 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoL2E_000 <- mkReg(unpack(0));

    rule count_fifoL2E_000;

        let x_0 = (countDone_fifoL2E_000);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoL2E_000);
        counter_fifoL2E_000 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoL2E_000);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoL2E_000);
            $display ("-- LR fifoL2E_000: %b %x %b %x %x %x %b %x %x %b %x %b %x %b %x", ((x_3).lr_ir_pp).ir_is_rs_rel, (((x_3).lr_ir_pp).ir_msg).id, (((x_3).lr_ir_pp).ir_msg).type_, (((x_3).lr_ir_pp).ir_msg).addr, ((x_3).lr_ir_pp).ir_msg_from, ((x_3).lr_ir_pp).ir_mshr_id, (((x_3).lr_ir_pp).ir_by_victim).valid, (((x_3).lr_ir_pp).ir_by_victim).data, ((x_3).lr_ir).info_index, ((x_3).lr_ir).info_hit, ((x_3).lr_ir).info_way, ((x_3).lr_ir).edir_hit, ((x_3).lr_ir).edir_way, (((x_3).lr_ir).edir_slot).valid, (((x_3).lr_ir).edir_slot).data);
            countDone_fifoL2E_000 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoL2E_000 (Struct43 x_0);
        let x_1 = (full_fifoL2E_000);
        when (! (x_1), noAction);
        elt_fifoL2E_000 <= x_0;
        full_fifoL2E_000 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct43) deq_fifoL2E_000 ();
        let x_1 = (full_fifoL2E_000);
        when (x_1, noAction);
        let x_2 = (elt_fifoL2E_000);
        full_fifoL2E_000 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module40;
    method Action enq_fifo0000 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0000 ();
endinterface

module mkModule40
    (Module40);
    Reg#(Vector#(2, Struct1)) elt_fifo0000 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0000 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0000 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0000 <- mkReg(True);
    Reg#(Bool) full_fifo0000 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0000 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0000 <- mkReg(unpack(0));

    rule count_fifo0000;

        let x_0 = (countDone_fifo0000);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0000);
        counter_fifo0000 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0000);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0000);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0000:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0000:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0000 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0000 (Struct1 x_0);
        let x_1 = (full_fifo0000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0000);
        let x_3 = (enqP_fifo0000);
        let x_4 = (deqP_fifo0000);
        elt_fifo0000 <= update (x_2, x_3, x_0);
        empty_fifo0000 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0000 <= (x_4) == (x_5);
        enqP_fifo0000 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0000 ();
        let x_1 = (empty_fifo0000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0000);
        let x_3 = (enqP_fifo0000);
        let x_4 = (deqP_fifo0000);
        full_fifo0000 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0000 <= (x_3) == (x_5);
        deqP_fifo0000 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module41;
    method Action enq_fifo0001 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0001 ();
endinterface

module mkModule41
    (Module41);
    Reg#(Vector#(2, Struct1)) elt_fifo0001 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0001 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0001 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0001 <- mkReg(True);
    Reg#(Bool) full_fifo0001 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0001 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0001 <- mkReg(unpack(0));

    rule count_fifo0001;

        let x_0 = (countDone_fifo0001);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0001);
        counter_fifo0001 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0001);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0001);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0001:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0001:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0001 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0001 (Struct1 x_0);
        let x_1 = (full_fifo0001);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0001);
        let x_3 = (enqP_fifo0001);
        let x_4 = (deqP_fifo0001);
        elt_fifo0001 <= update (x_2, x_3, x_0);
        empty_fifo0001 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0001 <= (x_4) == (x_5);
        enqP_fifo0001 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0001 ();
        let x_1 = (empty_fifo0001);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0001);
        let x_3 = (enqP_fifo0001);
        let x_4 = (deqP_fifo0001);
        full_fifo0001 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0001 <= (x_3) == (x_5);
        deqP_fifo0001 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module42;
    method Action enq_fifo0002 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0002 ();
endinterface

module mkModule42
    (Module42);
    Reg#(Vector#(2, Struct1)) elt_fifo0002 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0002 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0002 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0002 <- mkReg(True);
    Reg#(Bool) full_fifo0002 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0002 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0002 <- mkReg(unpack(0));

    rule count_fifo0002;

        let x_0 = (countDone_fifo0002);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0002);
        counter_fifo0002 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0002);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0002);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0002:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0002:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0002 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0002 (Struct1 x_0);
        let x_1 = (full_fifo0002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0002);
        let x_3 = (enqP_fifo0002);
        let x_4 = (deqP_fifo0002);
        elt_fifo0002 <= update (x_2, x_3, x_0);
        empty_fifo0002 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0002 <= (x_4) == (x_5);
        enqP_fifo0002 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0002 ();
        let x_1 = (empty_fifo0002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0002);
        let x_3 = (enqP_fifo0002);
        let x_4 = (deqP_fifo0002);
        full_fifo0002 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0002 <= (x_3) == (x_5);
        deqP_fifo0002 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module43;
    method Action enq_fifo00000 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00000 ();
endinterface

module mkModule43
    (Module43);
    Reg#(Vector#(2, Struct1)) elt_fifo00000 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00000 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00000 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00000 <- mkReg(True);
    Reg#(Bool) full_fifo00000 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00000 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00000 <- mkReg(unpack(0));

    rule count_fifo00000;

        let x_0 = (countDone_fifo00000);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00000);
        counter_fifo00000 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00000);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00000);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00000:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00000:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00000 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00000 (Struct1 x_0);
        let x_1 = (full_fifo00000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00000);
        let x_3 = (enqP_fifo00000);
        let x_4 = (deqP_fifo00000);
        elt_fifo00000 <= update (x_2, x_3, x_0);
        empty_fifo00000 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00000 <= (x_4) == (x_5);
        enqP_fifo00000 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00000 ();
        let x_1 = (empty_fifo00000);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00000);
        let x_3 = (enqP_fifo00000);
        let x_4 = (deqP_fifo00000);
        full_fifo00000 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00000 <= (x_3) == (x_5);
        deqP_fifo00000 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module44;
    method Action enq_fifo00002 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00002 ();
endinterface

module mkModule44
    (Module44);
    Reg#(Vector#(2, Struct1)) elt_fifo00002 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00002 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00002 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00002 <- mkReg(True);
    Reg#(Bool) full_fifo00002 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00002 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00002 <- mkReg(unpack(0));

    rule count_fifo00002;

        let x_0 = (countDone_fifo00002);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00002);
        counter_fifo00002 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00002);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00002);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00002:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00002:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00002 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00002 (Struct1 x_0);
        let x_1 = (full_fifo00002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00002);
        let x_3 = (enqP_fifo00002);
        let x_4 = (deqP_fifo00002);
        elt_fifo00002 <= update (x_2, x_3, x_0);
        empty_fifo00002 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00002 <= (x_4) == (x_5);
        enqP_fifo00002 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00002 ();
        let x_1 = (empty_fifo00002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00002);
        let x_3 = (enqP_fifo00002);
        let x_4 = (deqP_fifo00002);
        full_fifo00002 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00002 <= (x_3) == (x_5);
        deqP_fifo00002 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module45;
    method ActionValue#(Struct39) victims__000__findVictim (Bit#(64) x_0);
    method ActionValue#(Struct44) victims__000__getVictim (Bit#(2) x_0);
    method Action victims__000__setVictim (Struct48 x_0);
    method Action victims__000__registerVictim (Struct44 x_0);
    method ActionValue#(Struct44) victims__000__getFirstVictim ();
    method ActionValue#(Bool) victims__000__hasVictim ();
    method Action victims__000__setVictimRq (Struct49 x_0);
    method ActionValue#(Bit#(3)) victims__000__releaseVictim (Bit#(64) x_0);
endinterface

module mkModule45
    (Module45);
    Reg#(Vector#(4, Struct44)) victimRegs__000 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct39) victims__000__findVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__000);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_9 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            x_9 = Struct39 {valid : (Bool)'(True), data : (Bit#(2))'(2'h0)};
        end else begin
            Struct44 x_3 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_8 = ?;
            if (((x_3).victim_valid) && (((x_3).victim_addr) == (x_0)))
                begin
                x_8 = Struct39 {valid : (Bool)'(True), data :
                (Bit#(2))'(2'h1)};
            end else begin
                Struct44 x_4 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_7 = ?;
                if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                    begin
                    x_7 = Struct39 {valid : (Bool)'(True), data :
                    (Bit#(2))'(2'h2)};
                end else begin
                    Struct44 x_5 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_6 = ?;
                    if (((x_5).victim_valid) && (((x_5).victim_addr) ==
                        (x_0))) begin
                        x_6 = Struct39 {valid : (Bool)'(True), data :
                        (Bit#(2))'(2'h3)};
                    end else begin
                        x_6 = Struct39 {valid : (Bool)'(False), data :
                        unpack(0)};
                    end
                    x_7 = x_6;
                end
                x_8 = x_7;
            end
            x_9 = x_8;
        end
        return x_9;
    endmethod

    method ActionValue#(Struct44) victims__000__getVictim (Bit#(2) x_0);
        let x_1 = (victimRegs__000);
        return (x_1)[x_0];
    endmethod

    method Action victims__000__setVictim (Struct48 x_0);
        let x_1 = (victimRegs__000);
        Struct44 x_2 = ((x_1)[(x_0).victim_idx]);
        Struct44 x_3 = (Struct44 {victim_valid : (Bool)'(True), victim_addr :
        (x_2).victim_addr, victim_info : (x_0).victim_info, victim_value :
        (x_0).victim_value, victim_req : (x_2).victim_req});
        victimRegs__000 <= update (x_1, (x_0).victim_idx, x_3);
    endmethod

    method Action victims__000__registerVictim (Struct44 x_0);
        let x_1 = (victimRegs__000);
        Struct39 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_valid ? (Struct39 {valid :
        (Bool)'(False), data : unpack(0)}) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h0)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h1)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h2)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h3)})));
        when ((x_2).valid, noAction);
        Bit#(2) x_3 = ((x_2).data);
        victimRegs__000 <= update (x_1, x_3, x_0);
    endmethod

    method ActionValue#(Struct44) victims__000__getFirstVictim ();
        let x_1 = (victimRegs__000);
        Struct55 x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) : (Struct55 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method ActionValue#(Bool) victims__000__hasVictim ();
        let x_1 = (victimRegs__000);
        Bool x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        return x_2;
    endmethod

    method Action victims__000__setVictimRq (Struct49 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victimRegs__000);
        Struct44 x_4 =
        ((x_3)[(Bit#(2))'(2'h3)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct44 x_5 = (Struct44 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct5 {valid :
            (Bool)'(True), data : x_2}});
            victimRegs__000 <= update (x_3, (Bit#(2))'(2'h3), x_5);
        end else begin
            Struct44 x_6 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct44 x_7 = (Struct44 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct5 {valid : (Bool)'(True), data :
                x_2}});
                victimRegs__000 <= update (x_3, (Bit#(2))'(2'h2), x_7);
            end else begin
                Struct44 x_8 =
                ((x_3)[(Bit#(2))'(2'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct44 x_9 = (Struct44 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct5 {valid :
                    (Bool)'(True), data : x_2}});
                    victimRegs__000 <= update (x_3, (Bit#(2))'(2'h1), x_9);
                end else begin
                    Struct44 x_10 =
                    ((x_3)[(Bit#(2))'(2'h0)]);
                    if (((x_10).victim_valid) && (((x_10).victim_addr) ==
                        (x_1))) begin
                        Struct44 x_11 = (Struct44 {victim_valid :
                        (x_10).victim_valid, victim_addr :
                        (x_10).victim_addr, victim_info : (x_10).victim_info,
                        victim_value : (x_10).victim_value, victim_req :
                        Struct5 {valid : (Bool)'(True), data :
                        x_2}});
                        victimRegs__000 <= update (x_3, (Bit#(2))'(2'h0),
                        x_11);
                    end else begin

                    end
                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) victims__000__releaseVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__000);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victimRegs__000 <= update (x_1, (Bit#(2))'(2'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct44 x_4 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victimRegs__000 <= update (x_1, (Bit#(2))'(2'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct44 x_6 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victimRegs__000 <= update (x_1, (Bit#(2))'(2'h2),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct44 x_8 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victimRegs__000 <= update (x_1, (Bit#(2))'(2'h3),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod
endmodule

interface Module46;
    method Action rdReq_infoRam__000__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__000__3 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__000__3 ();
endinterface

module mkModule46 (Module46);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h7, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__3 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__000__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module47;
    method Action rdReq_infoRam__000__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__000__2 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__000__2 ();
endinterface

module mkModule47 (Module47);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h6, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__2 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__000__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module48;
    method Action rdReq_infoRam__000__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__000__1 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__000__1 ();
endinterface

module mkModule48 (Module48);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h5, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__1 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__000__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module49;
    method Action rdReq_infoRam__000__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__000__0 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__000__0 ();
endinterface

module mkModule49 (Module49);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h4, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__0 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__000__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module50;
    method Action rdReq_dataRam__000 (Bit#(10) x_0);
    method Action wrReq_dataRam__000 (Struct54 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__000 ();
endinterface

module mkModule50 (Module50);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__000 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__000 (Struct54 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__000 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module51;
    method Action rdReq_repRam__000 (Bit#(8) x_0);
    method Action wrReq_repRam__000 (Struct56 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__000 ();
endinterface

module mkModule51 (Module51);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h1, 8'h1, 8'h1, 8'h1);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__000 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__000 (Struct56 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__000 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module52;
    method ActionValue#(Struct45) getMSHR_000 (Bit#(3) x_0);
    method ActionValue#(Struct38) getPRqSlot_000 (Struct37 x_0);
    method ActionValue#(Struct38) getCRqSlot_000 (Struct37 x_0);
    method ActionValue#(Struct37) getWait_000 ();
    method Action registerUL_000 (Struct47 x_0);
    method Action registerDL_000 (Struct57 x_0);
    method Action canImm_000 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) setULImm_000 (Struct1 x_0);
    method Action transferUpDown_000 (Struct58 x_0);
    method Action addRs_000 (Struct7 x_0);
    method ActionValue#(Bit#(3)) getULReady_000 (Bit#(64) x_0);
    method ActionValue#(Struct59) getDLReady_000 ();
    method Action startRelease_000 (Bit#(3) x_0);
    method Action releaseMSHR_000 (Bit#(3) x_0);
endinterface

module mkModule52
    (Module52);
    Reg#(Vector#(6, Struct45)) rqs_000 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct45) getMSHR_000 (Bit#(3) x_0);
        let x_1 = (rqs_000);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct38) getPRqSlot_000 (Struct37 x_0);
        let x_1 = (rqs_000);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_8 = ((x_7).valid);
        Struct38 x_9 = (Struct38 {s_has_slot : (x_3) && (! (x_6)), s_conflict
        : x_8, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_10 = (update (x_1, x_4, Struct45 {m_status
            : (x_8 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_14 = ?;
            if (x_8) begin
                Bit#(3) x_11 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
                ((Bit#(3))'(3'h0)))) && (!
                ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h0)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h1)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h2)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h3)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h4)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
                Struct45 x_12 = ((x_1)[x_11]);
                Vector#(6, Struct45) x_13 = (update (x_10, x_11, Struct45
                {m_status : (x_12).m_status, m_next : (x_8 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_12).m_next)), m_is_ul :
                (x_12).m_is_ul, m_msg : (x_12).m_msg, m_qidx : (x_12).m_qidx,
                m_rsb : (x_12).m_rsb, m_dl_rss_from : (x_12).m_dl_rss_from,
                m_dl_rss_recv : (x_12).m_dl_rss_recv, m_dl_rss :
                (x_12).m_dl_rss}));
                x_14 = x_13;
            end else begin
                x_14 = x_10;
            end
            rqs_000 <= x_14;
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct38) getCRqSlot_000 (Struct37 x_0);
        let x_1 = (rqs_000);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        Struct5 x_8 = (((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_9 = ((x_7).valid);
        Bool x_10 = ((x_8).valid);
        Bool x_11 = ((x_9) || (x_10));
        Struct38 x_12 = (Struct38 {s_has_slot : (x_3) && (! (x_6)),
        s_conflict : x_11, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_13 = (update (x_1, x_4, Struct45 {m_status
            : (x_11 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_17 = ?;
            if (x_11) begin
                Bit#(3) x_14 = ((x_9 ? ((x_7).data) : ((x_8).data)));
                Struct45 x_15 = ((x_1)[x_14]);
                Vector#(6, Struct45) x_16 = (update (x_13, x_14, Struct45
                {m_status : (x_15).m_status, m_next : (x_11 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_15).m_next)), m_is_ul :
                (x_15).m_is_ul, m_msg : (x_15).m_msg, m_qidx : (x_15).m_qidx,
                m_rsb : (x_15).m_rsb, m_dl_rss_from : (x_15).m_dl_rss_from,
                m_dl_rss_recv : (x_15).m_dl_rss_recv, m_dl_rss :
                (x_15).m_dl_rss}));
                x_17 = x_16;
            end else begin
                x_17 = x_13;
            end
            rqs_000 <= x_17;
        end else begin

        end
        return x_12;
    endmethod

    method ActionValue#(Struct37) getWait_000 ();
        let x_1 = (rqs_000);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h4)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        rqs_000 <= update (x_1, x_3, Struct45 {m_status : (Bit#(3))'(3'h4),
        m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg,
        m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : (x_4).m_dl_rss_recv, m_dl_rss :
        (x_4).m_dl_rss});
        Struct37 x_7 = (Struct37 {r_id : x_3, r_msg : (x_4).m_msg, r_msg_from
        : (x_4).m_qidx});
        return x_7;
    endmethod

    method Action registerUL_000 (Struct47 x_0);
        let x_1 = (rqs_000);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_000 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_000 (Struct57 x_0);
        let x_1 = (rqs_000);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_000 <= update (x_1, x_2, x_4);
    endmethod

    method Action canImm_000 (Bit#(64) x_0);
        let x_1 = (rqs_000);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
    endmethod

    method ActionValue#(Bit#(3)) setULImm_000 (Struct1 x_0);
        let x_1 = (rqs_000);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Bit#(64) x_4 = ((x_0).addr);
        Struct5 x_5 = (((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_4)) ? (Struct5 {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((! ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_5).valid), noAction);
        Vector#(6, Struct45) x_6 = (update (x_1, x_3, Struct45 {m_status :
        (Bit#(3))'(3'h5), m_next : Struct5 {valid : (Bool)'(False), data :
        unpack(0)}, m_is_ul : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)}));
        rqs_000 <= x_6;
        return x_3;
    endmethod

    method Action transferUpDown_000 (Struct58 x_0);
        let x_1 = (rqs_000);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_000 <= update (x_1, x_2, x_4);
    endmethod

    method Action addRs_000 (Struct7 x_0);
        let x_1 = (rqs_000);
        Bit#(64) x_2 = (((x_0).r_msg).addr);
        Struct5 x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_3).valid, noAction);
        Bit#(3) x_4 = ((x_3).data);
        Struct45 x_5 = ((x_1)[x_4]);
        Struct45 x_6 = (Struct45 {m_status : (x_5).m_status, m_next :
        (x_5).m_next, m_is_ul : (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx :
        (x_5).m_qidx, m_rsb : (x_5).m_rsb, m_dl_rss_from :
        (x_5).m_dl_rss_from, m_dl_rss_recv : ((x_5).m_dl_rss_recv) |
        (((Bit#(4))'(4'h1)) << ((x_0).r_midx)), m_dl_rss : update
        ((x_5).m_dl_rss, (x_0).r_midx, (x_0).r_msg)});
        rqs_000 <= update (x_1, x_4, x_6);
    endmethod

    method ActionValue#(Bit#(3)) getULReady_000 (Bit#(64) x_0);
        let x_1 = (rqs_000);
        Bool x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_2), noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
        Struct5 x_4 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_4).valid, noAction);
        Bit#(3) x_5 = ((x_4).data);
        return x_5;
    endmethod

    method ActionValue#(Struct59) getDLReady_000 ();
        let x_1 = (rqs_000);
        Struct5 x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        Struct59 x_7 = (Struct59 {r_id : x_3, r_addr : x_5});
        return x_7;
    endmethod

    method Action startRelease_000 (Bit#(3) x_0);
        let x_1 = (rqs_000);
        Struct45 x_2 = ((x_1)[x_0]);
        Struct45 x_3 = (Struct45 {m_status : (Bit#(3))'(3'h6), m_next :
        (x_2).m_next, m_is_ul : (x_2).m_is_ul, m_msg : (x_2).m_msg, m_qidx :
        (x_2).m_qidx, m_rsb : (x_2).m_rsb, m_dl_rss_from :
        (x_2).m_dl_rss_from, m_dl_rss_recv : (x_2).m_dl_rss_recv, m_dl_rss :
        (x_2).m_dl_rss});
        rqs_000 <= update (x_1, x_0, x_3);
    endmethod

    method Action releaseMSHR_000 (Bit#(3) x_0);
        let x_1 = (rqs_000);
        Struct45 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct45) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct45 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct45) x_6 = (update (x_3, x_4, Struct45 {m_status
            : (Bit#(3))'(3'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_000 <= x_7;
    endmethod
endmodule

interface Module53;
    method Action enq_fifoCRqInput_001 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput_001 ();
endinterface

module mkModule53
    (Module53);
    Reg#(Vector#(4, Struct2)) elt_fifoCRqInput_001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoCRqInput_001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoCRqInput_001 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoCRqInput_001 <- mkReg(True);
    Reg#(Bool) full_fifoCRqInput_001 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoCRqInput_001 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoCRqInput_001 <- mkReg(unpack(0));

    rule count_fifoCRqInput_001;

        let x_0 = (countDone_fifoCRqInput_001);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoCRqInput_001);
        counter_fifoCRqInput_001 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoCRqInput_001);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoCRqInput_001);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoCRqInput_001:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoCRqInput_001:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoCRqInput_001:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoCRqInput_001:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoCRqInput_001 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoCRqInput_001 (Struct2 x_0);
        let x_1 = (full_fifoCRqInput_001);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_001);
        let x_3 = (enqP_fifoCRqInput_001);
        let x_4 = (deqP_fifoCRqInput_001);
        elt_fifoCRqInput_001 <= update (x_2, x_3, x_0);
        empty_fifoCRqInput_001 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoCRqInput_001 <= (x_4) == (x_5);
        enqP_fifoCRqInput_001 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput_001 ();
        let x_1 = (empty_fifoCRqInput_001);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_001);
        let x_3 = (enqP_fifoCRqInput_001);
        let x_4 = (deqP_fifoCRqInput_001);
        full_fifoCRqInput_001 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoCRqInput_001 <= (x_3) == (x_5);
        deqP_fifoCRqInput_001 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module54;
    method Action enq_fifoPInput_001 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoPInput_001 ();
endinterface

module mkModule54
    (Module54);
    Reg#(Vector#(4, Struct2)) elt_fifoPInput_001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoPInput_001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoPInput_001 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoPInput_001 <- mkReg(True);
    Reg#(Bool) full_fifoPInput_001 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoPInput_001 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoPInput_001 <- mkReg(unpack(0));

    rule count_fifoPInput_001;

        let x_0 = (countDone_fifoPInput_001);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoPInput_001);
        counter_fifoPInput_001 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoPInput_001);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoPInput_001);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoPInput_001:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoPInput_001:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoPInput_001:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoPInput_001:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoPInput_001 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoPInput_001 (Struct2 x_0);
        let x_1 = (full_fifoPInput_001);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_001);
        let x_3 = (enqP_fifoPInput_001);
        let x_4 = (deqP_fifoPInput_001);
        elt_fifoPInput_001 <= update (x_2, x_3, x_0);
        empty_fifoPInput_001 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoPInput_001 <= (x_4) == (x_5);
        enqP_fifoPInput_001 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoPInput_001 ();
        let x_1 = (empty_fifoPInput_001);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_001);
        let x_3 = (enqP_fifoPInput_001);
        let x_4 = (deqP_fifoPInput_001);
        full_fifoPInput_001 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoPInput_001 <= (x_3) == (x_5);
        deqP_fifoPInput_001 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module55;
    method Action enq_fifoN2I_001 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoN2I_001 ();
endinterface

module mkModule55
    (Module55);
    Reg#(Struct40) elt_fifoN2I_001 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoN2I_001 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoN2I_001 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoN2I_001 <- mkReg(unpack(0));

    rule count_fifoN2I_001;

        let x_0 = (countDone_fifoN2I_001);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoN2I_001);
        counter_fifoN2I_001 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoN2I_001);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoN2I_001);
            $display ("-- IR fifoN2I_001: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoN2I_001 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoN2I_001 (Struct40 x_0);
        let x_1 = (full_fifoN2I_001);
        when (! (x_1), noAction);
        elt_fifoN2I_001 <= x_0;
        full_fifoN2I_001 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoN2I_001 ();
        let x_1 = (full_fifoN2I_001);
        when (x_1, noAction);
        let x_2 = (elt_fifoN2I_001);
        full_fifoN2I_001 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module56;
    method Action enq_fifoI2L_001 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoI2L_001 ();
endinterface

module mkModule56
    (Module56);
    Reg#(Struct40) elt_fifoI2L_001 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoI2L_001 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoI2L_001 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoI2L_001 <- mkReg(unpack(0));

    rule count_fifoI2L_001;

        let x_0 = (countDone_fifoI2L_001);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoI2L_001);
        counter_fifoI2L_001 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoI2L_001);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoI2L_001);
            $display ("-- IR fifoI2L_001: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoI2L_001 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoI2L_001 (Struct40 x_0);
        let x_1 = (full_fifoI2L_001);
        when (! (x_1), noAction);
        elt_fifoI2L_001 <= x_0;
        full_fifoI2L_001 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoI2L_001 ();
        let x_1 = (full_fifoI2L_001);
        when (x_1, noAction);
        let x_2 = (elt_fifoI2L_001);
        full_fifoI2L_001 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module57;
    method Action enq_fifoL2E_001 (Struct43 x_0);
    method ActionValue#(Struct43) deq_fifoL2E_001 ();
endinterface

module mkModule57
    (Module57);
    Reg#(Struct43) elt_fifoL2E_001 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoL2E_001 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoL2E_001 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoL2E_001 <- mkReg(unpack(0));

    rule count_fifoL2E_001;

        let x_0 = (countDone_fifoL2E_001);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoL2E_001);
        counter_fifoL2E_001 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoL2E_001);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoL2E_001);
            $display ("-- LR fifoL2E_001: %b %x %b %x %x %x %b %x %x %b %x %b %x %b %x", ((x_3).lr_ir_pp).ir_is_rs_rel, (((x_3).lr_ir_pp).ir_msg).id, (((x_3).lr_ir_pp).ir_msg).type_, (((x_3).lr_ir_pp).ir_msg).addr, ((x_3).lr_ir_pp).ir_msg_from, ((x_3).lr_ir_pp).ir_mshr_id, (((x_3).lr_ir_pp).ir_by_victim).valid, (((x_3).lr_ir_pp).ir_by_victim).data, ((x_3).lr_ir).info_index, ((x_3).lr_ir).info_hit, ((x_3).lr_ir).info_way, ((x_3).lr_ir).edir_hit, ((x_3).lr_ir).edir_way, (((x_3).lr_ir).edir_slot).valid, (((x_3).lr_ir).edir_slot).data);
            countDone_fifoL2E_001 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoL2E_001 (Struct43 x_0);
        let x_1 = (full_fifoL2E_001);
        when (! (x_1), noAction);
        elt_fifoL2E_001 <= x_0;
        full_fifoL2E_001 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct43) deq_fifoL2E_001 ();
        let x_1 = (full_fifoL2E_001);
        when (x_1, noAction);
        let x_2 = (elt_fifoL2E_001);
        full_fifoL2E_001 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module58;
    method Action enq_fifo0010 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0010 ();
endinterface

module mkModule58
    (Module58);
    Reg#(Vector#(2, Struct1)) elt_fifo0010 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0010 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0010 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0010 <- mkReg(True);
    Reg#(Bool) full_fifo0010 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0010 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0010 <- mkReg(unpack(0));

    rule count_fifo0010;

        let x_0 = (countDone_fifo0010);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0010);
        counter_fifo0010 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0010);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0010);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0010:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0010:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0010 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0010 (Struct1 x_0);
        let x_1 = (full_fifo0010);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0010);
        let x_3 = (enqP_fifo0010);
        let x_4 = (deqP_fifo0010);
        elt_fifo0010 <= update (x_2, x_3, x_0);
        empty_fifo0010 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0010 <= (x_4) == (x_5);
        enqP_fifo0010 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0010 ();
        let x_1 = (empty_fifo0010);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0010);
        let x_3 = (enqP_fifo0010);
        let x_4 = (deqP_fifo0010);
        full_fifo0010 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0010 <= (x_3) == (x_5);
        deqP_fifo0010 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module59;
    method Action enq_fifo0011 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0011 ();
endinterface

module mkModule59
    (Module59);
    Reg#(Vector#(2, Struct1)) elt_fifo0011 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0011 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0011 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0011 <- mkReg(True);
    Reg#(Bool) full_fifo0011 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0011 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0011 <- mkReg(unpack(0));

    rule count_fifo0011;

        let x_0 = (countDone_fifo0011);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0011);
        counter_fifo0011 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0011);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0011);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0011:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0011:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0011 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0011 (Struct1 x_0);
        let x_1 = (full_fifo0011);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0011);
        let x_3 = (enqP_fifo0011);
        let x_4 = (deqP_fifo0011);
        elt_fifo0011 <= update (x_2, x_3, x_0);
        empty_fifo0011 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0011 <= (x_4) == (x_5);
        enqP_fifo0011 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0011 ();
        let x_1 = (empty_fifo0011);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0011);
        let x_3 = (enqP_fifo0011);
        let x_4 = (deqP_fifo0011);
        full_fifo0011 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0011 <= (x_3) == (x_5);
        deqP_fifo0011 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module60;
    method Action enq_fifo0012 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0012 ();
endinterface

module mkModule60
    (Module60);
    Reg#(Vector#(2, Struct1)) elt_fifo0012 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0012 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0012 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0012 <- mkReg(True);
    Reg#(Bool) full_fifo0012 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0012 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0012 <- mkReg(unpack(0));

    rule count_fifo0012;

        let x_0 = (countDone_fifo0012);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0012);
        counter_fifo0012 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0012);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0012);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0012:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0012:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0012 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0012 (Struct1 x_0);
        let x_1 = (full_fifo0012);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0012);
        let x_3 = (enqP_fifo0012);
        let x_4 = (deqP_fifo0012);
        elt_fifo0012 <= update (x_2, x_3, x_0);
        empty_fifo0012 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0012 <= (x_4) == (x_5);
        enqP_fifo0012 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0012 ();
        let x_1 = (empty_fifo0012);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0012);
        let x_3 = (enqP_fifo0012);
        let x_4 = (deqP_fifo0012);
        full_fifo0012 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0012 <= (x_3) == (x_5);
        deqP_fifo0012 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module61;
    method Action enq_fifo00100 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00100 ();
endinterface

module mkModule61
    (Module61);
    Reg#(Vector#(2, Struct1)) elt_fifo00100 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00100 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00100 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00100 <- mkReg(True);
    Reg#(Bool) full_fifo00100 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00100 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00100 <- mkReg(unpack(0));

    rule count_fifo00100;

        let x_0 = (countDone_fifo00100);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00100);
        counter_fifo00100 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00100);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00100);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00100:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00100:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00100 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00100 (Struct1 x_0);
        let x_1 = (full_fifo00100);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00100);
        let x_3 = (enqP_fifo00100);
        let x_4 = (deqP_fifo00100);
        elt_fifo00100 <= update (x_2, x_3, x_0);
        empty_fifo00100 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00100 <= (x_4) == (x_5);
        enqP_fifo00100 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00100 ();
        let x_1 = (empty_fifo00100);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00100);
        let x_3 = (enqP_fifo00100);
        let x_4 = (deqP_fifo00100);
        full_fifo00100 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00100 <= (x_3) == (x_5);
        deqP_fifo00100 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module62;
    method Action enq_fifo00102 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00102 ();
endinterface

module mkModule62
    (Module62);
    Reg#(Vector#(2, Struct1)) elt_fifo00102 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00102 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00102 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00102 <- mkReg(True);
    Reg#(Bool) full_fifo00102 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00102 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00102 <- mkReg(unpack(0));

    rule count_fifo00102;

        let x_0 = (countDone_fifo00102);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00102);
        counter_fifo00102 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00102);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00102);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00102:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00102:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00102 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00102 (Struct1 x_0);
        let x_1 = (full_fifo00102);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00102);
        let x_3 = (enqP_fifo00102);
        let x_4 = (deqP_fifo00102);
        elt_fifo00102 <= update (x_2, x_3, x_0);
        empty_fifo00102 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00102 <= (x_4) == (x_5);
        enqP_fifo00102 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00102 ();
        let x_1 = (empty_fifo00102);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00102);
        let x_3 = (enqP_fifo00102);
        let x_4 = (deqP_fifo00102);
        full_fifo00102 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00102 <= (x_3) == (x_5);
        deqP_fifo00102 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module63;
    method ActionValue#(Struct39) victims__001__findVictim (Bit#(64) x_0);
    method ActionValue#(Struct44) victims__001__getVictim (Bit#(2) x_0);
    method Action victims__001__setVictim (Struct48 x_0);
    method Action victims__001__registerVictim (Struct44 x_0);
    method ActionValue#(Struct44) victims__001__getFirstVictim ();
    method ActionValue#(Bool) victims__001__hasVictim ();
    method Action victims__001__setVictimRq (Struct49 x_0);
    method ActionValue#(Bit#(3)) victims__001__releaseVictim (Bit#(64) x_0);
endinterface

module mkModule63
    (Module63);
    Reg#(Vector#(4, Struct44)) victimRegs__001 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct39) victims__001__findVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__001);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_9 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            x_9 = Struct39 {valid : (Bool)'(True), data : (Bit#(2))'(2'h0)};
        end else begin
            Struct44 x_3 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_8 = ?;
            if (((x_3).victim_valid) && (((x_3).victim_addr) == (x_0)))
                begin
                x_8 = Struct39 {valid : (Bool)'(True), data :
                (Bit#(2))'(2'h1)};
            end else begin
                Struct44 x_4 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_7 = ?;
                if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                    begin
                    x_7 = Struct39 {valid : (Bool)'(True), data :
                    (Bit#(2))'(2'h2)};
                end else begin
                    Struct44 x_5 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_6 = ?;
                    if (((x_5).victim_valid) && (((x_5).victim_addr) ==
                        (x_0))) begin
                        x_6 = Struct39 {valid : (Bool)'(True), data :
                        (Bit#(2))'(2'h3)};
                    end else begin
                        x_6 = Struct39 {valid : (Bool)'(False), data :
                        unpack(0)};
                    end
                    x_7 = x_6;
                end
                x_8 = x_7;
            end
            x_9 = x_8;
        end
        return x_9;
    endmethod

    method ActionValue#(Struct44) victims__001__getVictim (Bit#(2) x_0);
        let x_1 = (victimRegs__001);
        return (x_1)[x_0];
    endmethod

    method Action victims__001__setVictim (Struct48 x_0);
        let x_1 = (victimRegs__001);
        Struct44 x_2 = ((x_1)[(x_0).victim_idx]);
        Struct44 x_3 = (Struct44 {victim_valid : (Bool)'(True), victim_addr :
        (x_2).victim_addr, victim_info : (x_0).victim_info, victim_value :
        (x_0).victim_value, victim_req : (x_2).victim_req});
        victimRegs__001 <= update (x_1, (x_0).victim_idx, x_3);
    endmethod

    method Action victims__001__registerVictim (Struct44 x_0);
        let x_1 = (victimRegs__001);
        Struct39 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_valid ? (Struct39 {valid :
        (Bool)'(False), data : unpack(0)}) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h0)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h1)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h2)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h3)})));
        when ((x_2).valid, noAction);
        Bit#(2) x_3 = ((x_2).data);
        victimRegs__001 <= update (x_1, x_3, x_0);
    endmethod

    method ActionValue#(Struct44) victims__001__getFirstVictim ();
        let x_1 = (victimRegs__001);
        Struct55 x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) : (Struct55 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method ActionValue#(Bool) victims__001__hasVictim ();
        let x_1 = (victimRegs__001);
        Bool x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        return x_2;
    endmethod

    method Action victims__001__setVictimRq (Struct49 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victimRegs__001);
        Struct44 x_4 =
        ((x_3)[(Bit#(2))'(2'h3)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct44 x_5 = (Struct44 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct5 {valid :
            (Bool)'(True), data : x_2}});
            victimRegs__001 <= update (x_3, (Bit#(2))'(2'h3), x_5);
        end else begin
            Struct44 x_6 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct44 x_7 = (Struct44 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct5 {valid : (Bool)'(True), data :
                x_2}});
                victimRegs__001 <= update (x_3, (Bit#(2))'(2'h2), x_7);
            end else begin
                Struct44 x_8 =
                ((x_3)[(Bit#(2))'(2'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct44 x_9 = (Struct44 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct5 {valid :
                    (Bool)'(True), data : x_2}});
                    victimRegs__001 <= update (x_3, (Bit#(2))'(2'h1), x_9);
                end else begin
                    Struct44 x_10 =
                    ((x_3)[(Bit#(2))'(2'h0)]);
                    if (((x_10).victim_valid) && (((x_10).victim_addr) ==
                        (x_1))) begin
                        Struct44 x_11 = (Struct44 {victim_valid :
                        (x_10).victim_valid, victim_addr :
                        (x_10).victim_addr, victim_info : (x_10).victim_info,
                        victim_value : (x_10).victim_value, victim_req :
                        Struct5 {valid : (Bool)'(True), data :
                        x_2}});
                        victimRegs__001 <= update (x_3, (Bit#(2))'(2'h0),
                        x_11);
                    end else begin

                    end
                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) victims__001__releaseVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__001);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victimRegs__001 <= update (x_1, (Bit#(2))'(2'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct44 x_4 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victimRegs__001 <= update (x_1, (Bit#(2))'(2'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct44 x_6 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victimRegs__001 <= update (x_1, (Bit#(2))'(2'h2),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct44 x_8 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victimRegs__001 <= update (x_1, (Bit#(2))'(2'h3),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod
endmodule

interface Module64;
    method Action rdReq_infoRam__001__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__001__3 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__001__3 ();
endinterface

module mkModule64 (Module64);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h7, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__3 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__001__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module65;
    method Action rdReq_infoRam__001__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__001__2 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__001__2 ();
endinterface

module mkModule65 (Module65);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h6, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__2 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__001__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module66;
    method Action rdReq_infoRam__001__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__001__1 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__001__1 ();
endinterface

module mkModule66 (Module66);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h5, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__1 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__001__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module67;
    method Action rdReq_infoRam__001__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__001__0 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__001__0 ();
endinterface

module mkModule67 (Module67);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h4, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__0 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__001__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module68;
    method Action rdReq_dataRam__001 (Bit#(10) x_0);
    method Action wrReq_dataRam__001 (Struct54 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__001 ();
endinterface

module mkModule68 (Module68);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__001 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__001 (Struct54 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__001 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module69;
    method Action rdReq_repRam__001 (Bit#(8) x_0);
    method Action wrReq_repRam__001 (Struct56 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__001 ();
endinterface

module mkModule69 (Module69);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h1, 8'h1, 8'h1, 8'h1);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__001 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__001 (Struct56 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__001 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module70;
    method ActionValue#(Struct45) getMSHR_001 (Bit#(3) x_0);
    method ActionValue#(Struct38) getPRqSlot_001 (Struct37 x_0);
    method ActionValue#(Struct38) getCRqSlot_001 (Struct37 x_0);
    method ActionValue#(Struct37) getWait_001 ();
    method Action registerUL_001 (Struct47 x_0);
    method Action registerDL_001 (Struct57 x_0);
    method Action canImm_001 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) setULImm_001 (Struct1 x_0);
    method Action transferUpDown_001 (Struct58 x_0);
    method Action addRs_001 (Struct7 x_0);
    method ActionValue#(Bit#(3)) getULReady_001 (Bit#(64) x_0);
    method ActionValue#(Struct59) getDLReady_001 ();
    method Action startRelease_001 (Bit#(3) x_0);
    method Action releaseMSHR_001 (Bit#(3) x_0);
endinterface

module mkModule70
    (Module70);
    Reg#(Vector#(6, Struct45)) rqs_001 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct45) getMSHR_001 (Bit#(3) x_0);
        let x_1 = (rqs_001);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct38) getPRqSlot_001 (Struct37 x_0);
        let x_1 = (rqs_001);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_8 = ((x_7).valid);
        Struct38 x_9 = (Struct38 {s_has_slot : (x_3) && (! (x_6)), s_conflict
        : x_8, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_10 = (update (x_1, x_4, Struct45 {m_status
            : (x_8 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_14 = ?;
            if (x_8) begin
                Bit#(3) x_11 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
                ((Bit#(3))'(3'h0)))) && (!
                ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h0)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h1)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h2)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h3)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h4)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
                Struct45 x_12 = ((x_1)[x_11]);
                Vector#(6, Struct45) x_13 = (update (x_10, x_11, Struct45
                {m_status : (x_12).m_status, m_next : (x_8 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_12).m_next)), m_is_ul :
                (x_12).m_is_ul, m_msg : (x_12).m_msg, m_qidx : (x_12).m_qidx,
                m_rsb : (x_12).m_rsb, m_dl_rss_from : (x_12).m_dl_rss_from,
                m_dl_rss_recv : (x_12).m_dl_rss_recv, m_dl_rss :
                (x_12).m_dl_rss}));
                x_14 = x_13;
            end else begin
                x_14 = x_10;
            end
            rqs_001 <= x_14;
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct38) getCRqSlot_001 (Struct37 x_0);
        let x_1 = (rqs_001);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        Struct5 x_8 = (((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_9 = ((x_7).valid);
        Bool x_10 = ((x_8).valid);
        Bool x_11 = ((x_9) || (x_10));
        Struct38 x_12 = (Struct38 {s_has_slot : (x_3) && (! (x_6)),
        s_conflict : x_11, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_13 = (update (x_1, x_4, Struct45 {m_status
            : (x_11 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_17 = ?;
            if (x_11) begin
                Bit#(3) x_14 = ((x_9 ? ((x_7).data) : ((x_8).data)));
                Struct45 x_15 = ((x_1)[x_14]);
                Vector#(6, Struct45) x_16 = (update (x_13, x_14, Struct45
                {m_status : (x_15).m_status, m_next : (x_11 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_15).m_next)), m_is_ul :
                (x_15).m_is_ul, m_msg : (x_15).m_msg, m_qidx : (x_15).m_qidx,
                m_rsb : (x_15).m_rsb, m_dl_rss_from : (x_15).m_dl_rss_from,
                m_dl_rss_recv : (x_15).m_dl_rss_recv, m_dl_rss :
                (x_15).m_dl_rss}));
                x_17 = x_16;
            end else begin
                x_17 = x_13;
            end
            rqs_001 <= x_17;
        end else begin

        end
        return x_12;
    endmethod

    method ActionValue#(Struct37) getWait_001 ();
        let x_1 = (rqs_001);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h4)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        rqs_001 <= update (x_1, x_3, Struct45 {m_status : (Bit#(3))'(3'h4),
        m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg,
        m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : (x_4).m_dl_rss_recv, m_dl_rss :
        (x_4).m_dl_rss});
        Struct37 x_7 = (Struct37 {r_id : x_3, r_msg : (x_4).m_msg, r_msg_from
        : (x_4).m_qidx});
        return x_7;
    endmethod

    method Action registerUL_001 (Struct47 x_0);
        let x_1 = (rqs_001);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_001 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_001 (Struct57 x_0);
        let x_1 = (rqs_001);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_001 <= update (x_1, x_2, x_4);
    endmethod

    method Action canImm_001 (Bit#(64) x_0);
        let x_1 = (rqs_001);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
    endmethod

    method ActionValue#(Bit#(3)) setULImm_001 (Struct1 x_0);
        let x_1 = (rqs_001);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Bit#(64) x_4 = ((x_0).addr);
        Struct5 x_5 = (((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_4)) ? (Struct5 {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((! ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_5).valid), noAction);
        Vector#(6, Struct45) x_6 = (update (x_1, x_3, Struct45 {m_status :
        (Bit#(3))'(3'h5), m_next : Struct5 {valid : (Bool)'(False), data :
        unpack(0)}, m_is_ul : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)}));
        rqs_001 <= x_6;
        return x_3;
    endmethod

    method Action transferUpDown_001 (Struct58 x_0);
        let x_1 = (rqs_001);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_001 <= update (x_1, x_2, x_4);
    endmethod

    method Action addRs_001 (Struct7 x_0);
        let x_1 = (rqs_001);
        Bit#(64) x_2 = (((x_0).r_msg).addr);
        Struct5 x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_3).valid, noAction);
        Bit#(3) x_4 = ((x_3).data);
        Struct45 x_5 = ((x_1)[x_4]);
        Struct45 x_6 = (Struct45 {m_status : (x_5).m_status, m_next :
        (x_5).m_next, m_is_ul : (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx :
        (x_5).m_qidx, m_rsb : (x_5).m_rsb, m_dl_rss_from :
        (x_5).m_dl_rss_from, m_dl_rss_recv : ((x_5).m_dl_rss_recv) |
        (((Bit#(4))'(4'h1)) << ((x_0).r_midx)), m_dl_rss : update
        ((x_5).m_dl_rss, (x_0).r_midx, (x_0).r_msg)});
        rqs_001 <= update (x_1, x_4, x_6);
    endmethod

    method ActionValue#(Bit#(3)) getULReady_001 (Bit#(64) x_0);
        let x_1 = (rqs_001);
        Bool x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_2), noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
        Struct5 x_4 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_4).valid, noAction);
        Bit#(3) x_5 = ((x_4).data);
        return x_5;
    endmethod

    method ActionValue#(Struct59) getDLReady_001 ();
        let x_1 = (rqs_001);
        Struct5 x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        Struct59 x_7 = (Struct59 {r_id : x_3, r_addr : x_5});
        return x_7;
    endmethod

    method Action startRelease_001 (Bit#(3) x_0);
        let x_1 = (rqs_001);
        Struct45 x_2 = ((x_1)[x_0]);
        Struct45 x_3 = (Struct45 {m_status : (Bit#(3))'(3'h6), m_next :
        (x_2).m_next, m_is_ul : (x_2).m_is_ul, m_msg : (x_2).m_msg, m_qidx :
        (x_2).m_qidx, m_rsb : (x_2).m_rsb, m_dl_rss_from :
        (x_2).m_dl_rss_from, m_dl_rss_recv : (x_2).m_dl_rss_recv, m_dl_rss :
        (x_2).m_dl_rss});
        rqs_001 <= update (x_1, x_0, x_3);
    endmethod

    method Action releaseMSHR_001 (Bit#(3) x_0);
        let x_1 = (rqs_001);
        Struct45 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct45) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct45 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct45) x_6 = (update (x_3, x_4, Struct45 {m_status
            : (Bit#(3))'(3'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_001 <= x_7;
    endmethod
endmodule

interface Module71;
    method Action enq_fifoCRqInput_002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput_002 ();
endinterface

module mkModule71
    (Module71);
    Reg#(Vector#(4, Struct2)) elt_fifoCRqInput_002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoCRqInput_002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoCRqInput_002 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoCRqInput_002 <- mkReg(True);
    Reg#(Bool) full_fifoCRqInput_002 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoCRqInput_002 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoCRqInput_002 <- mkReg(unpack(0));

    rule count_fifoCRqInput_002;

        let x_0 = (countDone_fifoCRqInput_002);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoCRqInput_002);
        counter_fifoCRqInput_002 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoCRqInput_002);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoCRqInput_002);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoCRqInput_002:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoCRqInput_002:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoCRqInput_002:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoCRqInput_002:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoCRqInput_002 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoCRqInput_002 (Struct2 x_0);
        let x_1 = (full_fifoCRqInput_002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_002);
        let x_3 = (enqP_fifoCRqInput_002);
        let x_4 = (deqP_fifoCRqInput_002);
        elt_fifoCRqInput_002 <= update (x_2, x_3, x_0);
        empty_fifoCRqInput_002 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoCRqInput_002 <= (x_4) == (x_5);
        enqP_fifoCRqInput_002 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput_002 ();
        let x_1 = (empty_fifoCRqInput_002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_002);
        let x_3 = (enqP_fifoCRqInput_002);
        let x_4 = (deqP_fifoCRqInput_002);
        full_fifoCRqInput_002 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoCRqInput_002 <= (x_3) == (x_5);
        deqP_fifoCRqInput_002 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module72;
    method Action enq_fifoPInput_002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoPInput_002 ();
endinterface

module mkModule72
    (Module72);
    Reg#(Vector#(4, Struct2)) elt_fifoPInput_002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoPInput_002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoPInput_002 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoPInput_002 <- mkReg(True);
    Reg#(Bool) full_fifoPInput_002 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoPInput_002 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoPInput_002 <- mkReg(unpack(0));

    rule count_fifoPInput_002;

        let x_0 = (countDone_fifoPInput_002);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoPInput_002);
        counter_fifoPInput_002 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoPInput_002);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoPInput_002);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoPInput_002:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoPInput_002:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoPInput_002:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoPInput_002:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoPInput_002 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoPInput_002 (Struct2 x_0);
        let x_1 = (full_fifoPInput_002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_002);
        let x_3 = (enqP_fifoPInput_002);
        let x_4 = (deqP_fifoPInput_002);
        elt_fifoPInput_002 <= update (x_2, x_3, x_0);
        empty_fifoPInput_002 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoPInput_002 <= (x_4) == (x_5);
        enqP_fifoPInput_002 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoPInput_002 ();
        let x_1 = (empty_fifoPInput_002);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_002);
        let x_3 = (enqP_fifoPInput_002);
        let x_4 = (deqP_fifoPInput_002);
        full_fifoPInput_002 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoPInput_002 <= (x_3) == (x_5);
        deqP_fifoPInput_002 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module73;
    method Action enq_fifoN2I_002 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoN2I_002 ();
endinterface

module mkModule73
    (Module73);
    Reg#(Struct40) elt_fifoN2I_002 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoN2I_002 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoN2I_002 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoN2I_002 <- mkReg(unpack(0));

    rule count_fifoN2I_002;

        let x_0 = (countDone_fifoN2I_002);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoN2I_002);
        counter_fifoN2I_002 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoN2I_002);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoN2I_002);
            $display ("-- IR fifoN2I_002: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoN2I_002 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoN2I_002 (Struct40 x_0);
        let x_1 = (full_fifoN2I_002);
        when (! (x_1), noAction);
        elt_fifoN2I_002 <= x_0;
        full_fifoN2I_002 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoN2I_002 ();
        let x_1 = (full_fifoN2I_002);
        when (x_1, noAction);
        let x_2 = (elt_fifoN2I_002);
        full_fifoN2I_002 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module74;
    method Action enq_fifoI2L_002 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoI2L_002 ();
endinterface

module mkModule74
    (Module74);
    Reg#(Struct40) elt_fifoI2L_002 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoI2L_002 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoI2L_002 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoI2L_002 <- mkReg(unpack(0));

    rule count_fifoI2L_002;

        let x_0 = (countDone_fifoI2L_002);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoI2L_002);
        counter_fifoI2L_002 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoI2L_002);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoI2L_002);
            $display ("-- IR fifoI2L_002: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoI2L_002 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoI2L_002 (Struct40 x_0);
        let x_1 = (full_fifoI2L_002);
        when (! (x_1), noAction);
        elt_fifoI2L_002 <= x_0;
        full_fifoI2L_002 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoI2L_002 ();
        let x_1 = (full_fifoI2L_002);
        when (x_1, noAction);
        let x_2 = (elt_fifoI2L_002);
        full_fifoI2L_002 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module75;
    method Action enq_fifoL2E_002 (Struct43 x_0);
    method ActionValue#(Struct43) deq_fifoL2E_002 ();
endinterface

module mkModule75
    (Module75);
    Reg#(Struct43) elt_fifoL2E_002 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoL2E_002 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoL2E_002 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoL2E_002 <- mkReg(unpack(0));

    rule count_fifoL2E_002;

        let x_0 = (countDone_fifoL2E_002);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoL2E_002);
        counter_fifoL2E_002 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoL2E_002);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoL2E_002);
            $display ("-- LR fifoL2E_002: %b %x %b %x %x %x %b %x %x %b %x %b %x %b %x", ((x_3).lr_ir_pp).ir_is_rs_rel, (((x_3).lr_ir_pp).ir_msg).id, (((x_3).lr_ir_pp).ir_msg).type_, (((x_3).lr_ir_pp).ir_msg).addr, ((x_3).lr_ir_pp).ir_msg_from, ((x_3).lr_ir_pp).ir_mshr_id, (((x_3).lr_ir_pp).ir_by_victim).valid, (((x_3).lr_ir_pp).ir_by_victim).data, ((x_3).lr_ir).info_index, ((x_3).lr_ir).info_hit, ((x_3).lr_ir).info_way, ((x_3).lr_ir).edir_hit, ((x_3).lr_ir).edir_way, (((x_3).lr_ir).edir_slot).valid, (((x_3).lr_ir).edir_slot).data);
            countDone_fifoL2E_002 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoL2E_002 (Struct43 x_0);
        let x_1 = (full_fifoL2E_002);
        when (! (x_1), noAction);
        elt_fifoL2E_002 <= x_0;
        full_fifoL2E_002 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct43) deq_fifoL2E_002 ();
        let x_1 = (full_fifoL2E_002);
        when (x_1, noAction);
        let x_2 = (elt_fifoL2E_002);
        full_fifoL2E_002 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module76;
    method Action enq_fifo0020 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0020 ();
endinterface

module mkModule76
    (Module76);
    Reg#(Vector#(2, Struct1)) elt_fifo0020 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0020 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0020 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0020 <- mkReg(True);
    Reg#(Bool) full_fifo0020 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0020 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0020 <- mkReg(unpack(0));

    rule count_fifo0020;

        let x_0 = (countDone_fifo0020);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0020);
        counter_fifo0020 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0020);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0020);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0020:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0020:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0020 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0020 (Struct1 x_0);
        let x_1 = (full_fifo0020);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0020);
        let x_3 = (enqP_fifo0020);
        let x_4 = (deqP_fifo0020);
        elt_fifo0020 <= update (x_2, x_3, x_0);
        empty_fifo0020 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0020 <= (x_4) == (x_5);
        enqP_fifo0020 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0020 ();
        let x_1 = (empty_fifo0020);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0020);
        let x_3 = (enqP_fifo0020);
        let x_4 = (deqP_fifo0020);
        full_fifo0020 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0020 <= (x_3) == (x_5);
        deqP_fifo0020 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module77;
    method Action enq_fifo0021 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0021 ();
endinterface

module mkModule77
    (Module77);
    Reg#(Vector#(2, Struct1)) elt_fifo0021 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0021 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0021 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0021 <- mkReg(True);
    Reg#(Bool) full_fifo0021 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0021 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0021 <- mkReg(unpack(0));

    rule count_fifo0021;

        let x_0 = (countDone_fifo0021);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0021);
        counter_fifo0021 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0021);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0021);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0021:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0021:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0021 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0021 (Struct1 x_0);
        let x_1 = (full_fifo0021);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0021);
        let x_3 = (enqP_fifo0021);
        let x_4 = (deqP_fifo0021);
        elt_fifo0021 <= update (x_2, x_3, x_0);
        empty_fifo0021 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0021 <= (x_4) == (x_5);
        enqP_fifo0021 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0021 ();
        let x_1 = (empty_fifo0021);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0021);
        let x_3 = (enqP_fifo0021);
        let x_4 = (deqP_fifo0021);
        full_fifo0021 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0021 <= (x_3) == (x_5);
        deqP_fifo0021 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module78;
    method Action enq_fifo0022 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0022 ();
endinterface

module mkModule78
    (Module78);
    Reg#(Vector#(2, Struct1)) elt_fifo0022 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0022 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0022 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0022 <- mkReg(True);
    Reg#(Bool) full_fifo0022 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0022 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0022 <- mkReg(unpack(0));

    rule count_fifo0022;

        let x_0 = (countDone_fifo0022);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0022);
        counter_fifo0022 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0022);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0022);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0022:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0022:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0022 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0022 (Struct1 x_0);
        let x_1 = (full_fifo0022);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0022);
        let x_3 = (enqP_fifo0022);
        let x_4 = (deqP_fifo0022);
        elt_fifo0022 <= update (x_2, x_3, x_0);
        empty_fifo0022 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0022 <= (x_4) == (x_5);
        enqP_fifo0022 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0022 ();
        let x_1 = (empty_fifo0022);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0022);
        let x_3 = (enqP_fifo0022);
        let x_4 = (deqP_fifo0022);
        full_fifo0022 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0022 <= (x_3) == (x_5);
        deqP_fifo0022 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module79;
    method Action enq_fifo00200 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00200 ();
endinterface

module mkModule79
    (Module79);
    Reg#(Vector#(2, Struct1)) elt_fifo00200 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00200 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00200 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00200 <- mkReg(True);
    Reg#(Bool) full_fifo00200 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00200 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00200 <- mkReg(unpack(0));

    rule count_fifo00200;

        let x_0 = (countDone_fifo00200);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00200);
        counter_fifo00200 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00200);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00200);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00200:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00200:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00200 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00200 (Struct1 x_0);
        let x_1 = (full_fifo00200);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00200);
        let x_3 = (enqP_fifo00200);
        let x_4 = (deqP_fifo00200);
        elt_fifo00200 <= update (x_2, x_3, x_0);
        empty_fifo00200 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00200 <= (x_4) == (x_5);
        enqP_fifo00200 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00200 ();
        let x_1 = (empty_fifo00200);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00200);
        let x_3 = (enqP_fifo00200);
        let x_4 = (deqP_fifo00200);
        full_fifo00200 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00200 <= (x_3) == (x_5);
        deqP_fifo00200 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module80;
    method Action enq_fifo00202 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00202 ();
endinterface

module mkModule80
    (Module80);
    Reg#(Vector#(2, Struct1)) elt_fifo00202 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00202 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00202 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00202 <- mkReg(True);
    Reg#(Bool) full_fifo00202 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00202 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00202 <- mkReg(unpack(0));

    rule count_fifo00202;

        let x_0 = (countDone_fifo00202);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00202);
        counter_fifo00202 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00202);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00202);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00202:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00202:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00202 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00202 (Struct1 x_0);
        let x_1 = (full_fifo00202);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00202);
        let x_3 = (enqP_fifo00202);
        let x_4 = (deqP_fifo00202);
        elt_fifo00202 <= update (x_2, x_3, x_0);
        empty_fifo00202 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00202 <= (x_4) == (x_5);
        enqP_fifo00202 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00202 ();
        let x_1 = (empty_fifo00202);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00202);
        let x_3 = (enqP_fifo00202);
        let x_4 = (deqP_fifo00202);
        full_fifo00202 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00202 <= (x_3) == (x_5);
        deqP_fifo00202 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module81;
    method ActionValue#(Struct39) victims__002__findVictim (Bit#(64) x_0);
    method ActionValue#(Struct44) victims__002__getVictim (Bit#(2) x_0);
    method Action victims__002__setVictim (Struct48 x_0);
    method Action victims__002__registerVictim (Struct44 x_0);
    method ActionValue#(Struct44) victims__002__getFirstVictim ();
    method ActionValue#(Bool) victims__002__hasVictim ();
    method Action victims__002__setVictimRq (Struct49 x_0);
    method ActionValue#(Bit#(3)) victims__002__releaseVictim (Bit#(64) x_0);
endinterface

module mkModule81
    (Module81);
    Reg#(Vector#(4, Struct44)) victimRegs__002 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct39) victims__002__findVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__002);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_9 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            x_9 = Struct39 {valid : (Bool)'(True), data : (Bit#(2))'(2'h0)};
        end else begin
            Struct44 x_3 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_8 = ?;
            if (((x_3).victim_valid) && (((x_3).victim_addr) == (x_0)))
                begin
                x_8 = Struct39 {valid : (Bool)'(True), data :
                (Bit#(2))'(2'h1)};
            end else begin
                Struct44 x_4 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_7 = ?;
                if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                    begin
                    x_7 = Struct39 {valid : (Bool)'(True), data :
                    (Bit#(2))'(2'h2)};
                end else begin
                    Struct44 x_5 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_6 = ?;
                    if (((x_5).victim_valid) && (((x_5).victim_addr) ==
                        (x_0))) begin
                        x_6 = Struct39 {valid : (Bool)'(True), data :
                        (Bit#(2))'(2'h3)};
                    end else begin
                        x_6 = Struct39 {valid : (Bool)'(False), data :
                        unpack(0)};
                    end
                    x_7 = x_6;
                end
                x_8 = x_7;
            end
            x_9 = x_8;
        end
        return x_9;
    endmethod

    method ActionValue#(Struct44) victims__002__getVictim (Bit#(2) x_0);
        let x_1 = (victimRegs__002);
        return (x_1)[x_0];
    endmethod

    method Action victims__002__setVictim (Struct48 x_0);
        let x_1 = (victimRegs__002);
        Struct44 x_2 = ((x_1)[(x_0).victim_idx]);
        Struct44 x_3 = (Struct44 {victim_valid : (Bool)'(True), victim_addr :
        (x_2).victim_addr, victim_info : (x_0).victim_info, victim_value :
        (x_0).victim_value, victim_req : (x_2).victim_req});
        victimRegs__002 <= update (x_1, (x_0).victim_idx, x_3);
    endmethod

    method Action victims__002__registerVictim (Struct44 x_0);
        let x_1 = (victimRegs__002);
        Struct39 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_valid ? (Struct39 {valid :
        (Bool)'(False), data : unpack(0)}) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h0)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h1)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h2)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h3)})));
        when ((x_2).valid, noAction);
        Bit#(2) x_3 = ((x_2).data);
        victimRegs__002 <= update (x_1, x_3, x_0);
    endmethod

    method ActionValue#(Struct44) victims__002__getFirstVictim ();
        let x_1 = (victimRegs__002);
        Struct55 x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) : (Struct55 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method ActionValue#(Bool) victims__002__hasVictim ();
        let x_1 = (victimRegs__002);
        Bool x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        return x_2;
    endmethod

    method Action victims__002__setVictimRq (Struct49 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victimRegs__002);
        Struct44 x_4 =
        ((x_3)[(Bit#(2))'(2'h3)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct44 x_5 = (Struct44 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct5 {valid :
            (Bool)'(True), data : x_2}});
            victimRegs__002 <= update (x_3, (Bit#(2))'(2'h3), x_5);
        end else begin
            Struct44 x_6 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct44 x_7 = (Struct44 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct5 {valid : (Bool)'(True), data :
                x_2}});
                victimRegs__002 <= update (x_3, (Bit#(2))'(2'h2), x_7);
            end else begin
                Struct44 x_8 =
                ((x_3)[(Bit#(2))'(2'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct44 x_9 = (Struct44 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct5 {valid :
                    (Bool)'(True), data : x_2}});
                    victimRegs__002 <= update (x_3, (Bit#(2))'(2'h1), x_9);
                end else begin
                    Struct44 x_10 =
                    ((x_3)[(Bit#(2))'(2'h0)]);
                    if (((x_10).victim_valid) && (((x_10).victim_addr) ==
                        (x_1))) begin
                        Struct44 x_11 = (Struct44 {victim_valid :
                        (x_10).victim_valid, victim_addr :
                        (x_10).victim_addr, victim_info : (x_10).victim_info,
                        victim_value : (x_10).victim_value, victim_req :
                        Struct5 {valid : (Bool)'(True), data :
                        x_2}});
                        victimRegs__002 <= update (x_3, (Bit#(2))'(2'h0),
                        x_11);
                    end else begin

                    end
                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) victims__002__releaseVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__002);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victimRegs__002 <= update (x_1, (Bit#(2))'(2'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct44 x_4 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victimRegs__002 <= update (x_1, (Bit#(2))'(2'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct44 x_6 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victimRegs__002 <= update (x_1, (Bit#(2))'(2'h2),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct44 x_8 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victimRegs__002 <= update (x_1, (Bit#(2))'(2'h3),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod
endmodule

interface Module82;
    method Action rdReq_infoRam__002__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__002__3 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__002__3 ();
endinterface

module mkModule82 (Module82);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h7, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__002__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__002__3 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__002__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module83;
    method Action rdReq_infoRam__002__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__002__2 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__002__2 ();
endinterface

module mkModule83 (Module83);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h6, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__002__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__002__2 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__002__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module84;
    method Action rdReq_infoRam__002__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__002__1 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__002__1 ();
endinterface

module mkModule84 (Module84);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h5, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__002__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__002__1 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__002__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module85;
    method Action rdReq_infoRam__002__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__002__0 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__002__0 ();
endinterface

module mkModule85 (Module85);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h4, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__002__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__002__0 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__002__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module86;
    method Action rdReq_dataRam__002 (Bit#(10) x_0);
    method Action wrReq_dataRam__002 (Struct54 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__002 ();
endinterface

module mkModule86 (Module86);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__002 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__002 (Struct54 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__002 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module87;
    method Action rdReq_repRam__002 (Bit#(8) x_0);
    method Action wrReq_repRam__002 (Struct56 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__002 ();
endinterface

module mkModule87 (Module87);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h1, 8'h1, 8'h1, 8'h1);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__002 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__002 (Struct56 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__002 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module88;
    method ActionValue#(Struct45) getMSHR_002 (Bit#(3) x_0);
    method ActionValue#(Struct38) getPRqSlot_002 (Struct37 x_0);
    method ActionValue#(Struct38) getCRqSlot_002 (Struct37 x_0);
    method ActionValue#(Struct37) getWait_002 ();
    method Action registerUL_002 (Struct47 x_0);
    method Action registerDL_002 (Struct57 x_0);
    method Action canImm_002 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) setULImm_002 (Struct1 x_0);
    method Action transferUpDown_002 (Struct58 x_0);
    method Action addRs_002 (Struct7 x_0);
    method ActionValue#(Bit#(3)) getULReady_002 (Bit#(64) x_0);
    method ActionValue#(Struct59) getDLReady_002 ();
    method Action startRelease_002 (Bit#(3) x_0);
    method Action releaseMSHR_002 (Bit#(3) x_0);
endinterface

module mkModule88
    (Module88);
    Reg#(Vector#(6, Struct45)) rqs_002 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct45) getMSHR_002 (Bit#(3) x_0);
        let x_1 = (rqs_002);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct38) getPRqSlot_002 (Struct37 x_0);
        let x_1 = (rqs_002);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_8 = ((x_7).valid);
        Struct38 x_9 = (Struct38 {s_has_slot : (x_3) && (! (x_6)), s_conflict
        : x_8, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_10 = (update (x_1, x_4, Struct45 {m_status
            : (x_8 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_14 = ?;
            if (x_8) begin
                Bit#(3) x_11 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
                ((Bit#(3))'(3'h0)))) && (!
                ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h0)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h1)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h2)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h3)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h4)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
                Struct45 x_12 = ((x_1)[x_11]);
                Vector#(6, Struct45) x_13 = (update (x_10, x_11, Struct45
                {m_status : (x_12).m_status, m_next : (x_8 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_12).m_next)), m_is_ul :
                (x_12).m_is_ul, m_msg : (x_12).m_msg, m_qidx : (x_12).m_qidx,
                m_rsb : (x_12).m_rsb, m_dl_rss_from : (x_12).m_dl_rss_from,
                m_dl_rss_recv : (x_12).m_dl_rss_recv, m_dl_rss :
                (x_12).m_dl_rss}));
                x_14 = x_13;
            end else begin
                x_14 = x_10;
            end
            rqs_002 <= x_14;
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct38) getCRqSlot_002 (Struct37 x_0);
        let x_1 = (rqs_002);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        Struct5 x_8 = (((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_9 = ((x_7).valid);
        Bool x_10 = ((x_8).valid);
        Bool x_11 = ((x_9) || (x_10));
        Struct38 x_12 = (Struct38 {s_has_slot : (x_3) && (! (x_6)),
        s_conflict : x_11, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_13 = (update (x_1, x_4, Struct45 {m_status
            : (x_11 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_17 = ?;
            if (x_11) begin
                Bit#(3) x_14 = ((x_9 ? ((x_7).data) : ((x_8).data)));
                Struct45 x_15 = ((x_1)[x_14]);
                Vector#(6, Struct45) x_16 = (update (x_13, x_14, Struct45
                {m_status : (x_15).m_status, m_next : (x_11 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_15).m_next)), m_is_ul :
                (x_15).m_is_ul, m_msg : (x_15).m_msg, m_qidx : (x_15).m_qidx,
                m_rsb : (x_15).m_rsb, m_dl_rss_from : (x_15).m_dl_rss_from,
                m_dl_rss_recv : (x_15).m_dl_rss_recv, m_dl_rss :
                (x_15).m_dl_rss}));
                x_17 = x_16;
            end else begin
                x_17 = x_13;
            end
            rqs_002 <= x_17;
        end else begin

        end
        return x_12;
    endmethod

    method ActionValue#(Struct37) getWait_002 ();
        let x_1 = (rqs_002);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h4)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        rqs_002 <= update (x_1, x_3, Struct45 {m_status : (Bit#(3))'(3'h4),
        m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg,
        m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : (x_4).m_dl_rss_recv, m_dl_rss :
        (x_4).m_dl_rss});
        Struct37 x_7 = (Struct37 {r_id : x_3, r_msg : (x_4).m_msg, r_msg_from
        : (x_4).m_qidx});
        return x_7;
    endmethod

    method Action registerUL_002 (Struct47 x_0);
        let x_1 = (rqs_002);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_002 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_002 (Struct57 x_0);
        let x_1 = (rqs_002);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_002 <= update (x_1, x_2, x_4);
    endmethod

    method Action canImm_002 (Bit#(64) x_0);
        let x_1 = (rqs_002);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
    endmethod

    method ActionValue#(Bit#(3)) setULImm_002 (Struct1 x_0);
        let x_1 = (rqs_002);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Bit#(64) x_4 = ((x_0).addr);
        Struct5 x_5 = (((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_4)) ? (Struct5 {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((! ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_5).valid), noAction);
        Vector#(6, Struct45) x_6 = (update (x_1, x_3, Struct45 {m_status :
        (Bit#(3))'(3'h5), m_next : Struct5 {valid : (Bool)'(False), data :
        unpack(0)}, m_is_ul : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)}));
        rqs_002 <= x_6;
        return x_3;
    endmethod

    method Action transferUpDown_002 (Struct58 x_0);
        let x_1 = (rqs_002);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_002 <= update (x_1, x_2, x_4);
    endmethod

    method Action addRs_002 (Struct7 x_0);
        let x_1 = (rqs_002);
        Bit#(64) x_2 = (((x_0).r_msg).addr);
        Struct5 x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_3).valid, noAction);
        Bit#(3) x_4 = ((x_3).data);
        Struct45 x_5 = ((x_1)[x_4]);
        Struct45 x_6 = (Struct45 {m_status : (x_5).m_status, m_next :
        (x_5).m_next, m_is_ul : (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx :
        (x_5).m_qidx, m_rsb : (x_5).m_rsb, m_dl_rss_from :
        (x_5).m_dl_rss_from, m_dl_rss_recv : ((x_5).m_dl_rss_recv) |
        (((Bit#(4))'(4'h1)) << ((x_0).r_midx)), m_dl_rss : update
        ((x_5).m_dl_rss, (x_0).r_midx, (x_0).r_msg)});
        rqs_002 <= update (x_1, x_4, x_6);
    endmethod

    method ActionValue#(Bit#(3)) getULReady_002 (Bit#(64) x_0);
        let x_1 = (rqs_002);
        Bool x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_2), noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
        Struct5 x_4 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_4).valid, noAction);
        Bit#(3) x_5 = ((x_4).data);
        return x_5;
    endmethod

    method ActionValue#(Struct59) getDLReady_002 ();
        let x_1 = (rqs_002);
        Struct5 x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        Struct59 x_7 = (Struct59 {r_id : x_3, r_addr : x_5});
        return x_7;
    endmethod

    method Action startRelease_002 (Bit#(3) x_0);
        let x_1 = (rqs_002);
        Struct45 x_2 = ((x_1)[x_0]);
        Struct45 x_3 = (Struct45 {m_status : (Bit#(3))'(3'h6), m_next :
        (x_2).m_next, m_is_ul : (x_2).m_is_ul, m_msg : (x_2).m_msg, m_qidx :
        (x_2).m_qidx, m_rsb : (x_2).m_rsb, m_dl_rss_from :
        (x_2).m_dl_rss_from, m_dl_rss_recv : (x_2).m_dl_rss_recv, m_dl_rss :
        (x_2).m_dl_rss});
        rqs_002 <= update (x_1, x_0, x_3);
    endmethod

    method Action releaseMSHR_002 (Bit#(3) x_0);
        let x_1 = (rqs_002);
        Struct45 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct45) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct45 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct45) x_6 = (update (x_3, x_4, Struct45 {m_status
            : (Bit#(3))'(3'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_002 <= x_7;
    endmethod
endmodule

interface Module89;
    method Action enq_fifoCRqInput_003 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput_003 ();
endinterface

module mkModule89
    (Module89);
    Reg#(Vector#(4, Struct2)) elt_fifoCRqInput_003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoCRqInput_003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoCRqInput_003 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoCRqInput_003 <- mkReg(True);
    Reg#(Bool) full_fifoCRqInput_003 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoCRqInput_003 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoCRqInput_003 <- mkReg(unpack(0));

    rule count_fifoCRqInput_003;

        let x_0 = (countDone_fifoCRqInput_003);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoCRqInput_003);
        counter_fifoCRqInput_003 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoCRqInput_003);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoCRqInput_003);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoCRqInput_003:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoCRqInput_003:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoCRqInput_003:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoCRqInput_003:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoCRqInput_003 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoCRqInput_003 (Struct2 x_0);
        let x_1 = (full_fifoCRqInput_003);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_003);
        let x_3 = (enqP_fifoCRqInput_003);
        let x_4 = (deqP_fifoCRqInput_003);
        elt_fifoCRqInput_003 <= update (x_2, x_3, x_0);
        empty_fifoCRqInput_003 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoCRqInput_003 <= (x_4) == (x_5);
        enqP_fifoCRqInput_003 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput_003 ();
        let x_1 = (empty_fifoCRqInput_003);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoCRqInput_003);
        let x_3 = (enqP_fifoCRqInput_003);
        let x_4 = (deqP_fifoCRqInput_003);
        full_fifoCRqInput_003 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoCRqInput_003 <= (x_3) == (x_5);
        deqP_fifoCRqInput_003 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module90;
    method Action enq_fifoPInput_003 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoPInput_003 ();
endinterface

module mkModule90
    (Module90);
    Reg#(Vector#(4, Struct2)) elt_fifoPInput_003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) enqP_fifoPInput_003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) deqP_fifoPInput_003 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifoPInput_003 <- mkReg(True);
    Reg#(Bool) full_fifoPInput_003 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoPInput_003 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoPInput_003 <- mkReg(unpack(0));

    rule count_fifoPInput_003;

        let x_0 = (countDone_fifoPInput_003);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoPInput_003);
        counter_fifoPInput_003 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoPInput_003);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifoPInput_003);
            Struct2 x_4 =
            ((x_3)[(Bit#(2))'(2'h3)]);
            $display ("-- INPUT fifoPInput_003:3 %x %x %b %x", (x_4).in_msg_from, ((x_4).in_msg).id, ((x_4).in_msg).type_, ((x_4).in_msg).addr);
            Struct2 x_5 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            $display ("-- INPUT fifoPInput_003:2 %x %x %b %x", (x_5).in_msg_from, ((x_5).in_msg).id, ((x_5).in_msg).type_, ((x_5).in_msg).addr);
            Struct2 x_6 =
            ((x_3)[(Bit#(2))'(2'h1)]);
            $display ("-- INPUT fifoPInput_003:1 %x %x %b %x", (x_6).in_msg_from, ((x_6).in_msg).id, ((x_6).in_msg).type_, ((x_6).in_msg).addr);
            Struct2 x_7 =
            ((x_3)[(Bit#(2))'(2'h0)]);
            $display ("-- INPUT fifoPInput_003:0 %x %x %b %x", (x_7).in_msg_from, ((x_7).in_msg).id, ((x_7).in_msg).type_, ((x_7).in_msg).addr);
            countDone_fifoPInput_003 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoPInput_003 (Struct2 x_0);
        let x_1 = (full_fifoPInput_003);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_003);
        let x_3 = (enqP_fifoPInput_003);
        let x_4 = (deqP_fifoPInput_003);
        elt_fifoPInput_003 <= update (x_2, x_3, x_0);
        empty_fifoPInput_003 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_3) + ((Bit#(2))'(2'h1)));
        full_fifoPInput_003 <= (x_4) == (x_5);
        enqP_fifoPInput_003 <= x_5;
    endmethod

    method ActionValue#(Struct2) deq_fifoPInput_003 ();
        let x_1 = (empty_fifoPInput_003);
        when (! (x_1), noAction);
        let x_2 = (elt_fifoPInput_003);
        let x_3 = (enqP_fifoPInput_003);
        let x_4 = (deqP_fifoPInput_003);
        full_fifoPInput_003 <= (Bool)'(False);
        Bit#(2) x_5 = ((x_4) + ((Bit#(2))'(2'h1)));
        empty_fifoPInput_003 <= (x_3) == (x_5);
        deqP_fifoPInput_003 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module91;
    method Action enq_fifoN2I_003 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoN2I_003 ();
endinterface

module mkModule91
    (Module91);
    Reg#(Struct40) elt_fifoN2I_003 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoN2I_003 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoN2I_003 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoN2I_003 <- mkReg(unpack(0));

    rule count_fifoN2I_003;

        let x_0 = (countDone_fifoN2I_003);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoN2I_003);
        counter_fifoN2I_003 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoN2I_003);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoN2I_003);
            $display ("-- IR fifoN2I_003: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoN2I_003 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoN2I_003 (Struct40 x_0);
        let x_1 = (full_fifoN2I_003);
        when (! (x_1), noAction);
        elt_fifoN2I_003 <= x_0;
        full_fifoN2I_003 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoN2I_003 ();
        let x_1 = (full_fifoN2I_003);
        when (x_1, noAction);
        let x_2 = (elt_fifoN2I_003);
        full_fifoN2I_003 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module92;
    method Action enq_fifoI2L_003 (Struct40 x_0);
    method ActionValue#(Struct40) deq_fifoI2L_003 ();
endinterface

module mkModule92
    (Module92);
    Reg#(Struct40) elt_fifoI2L_003 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoI2L_003 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoI2L_003 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoI2L_003 <- mkReg(unpack(0));

    rule count_fifoI2L_003;

        let x_0 = (countDone_fifoI2L_003);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoI2L_003);
        counter_fifoI2L_003 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoI2L_003);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoI2L_003);
            $display ("-- IR fifoI2L_003: %b %x %b %x %x %x %b %x", (x_3).ir_is_rs_rel, ((x_3).ir_msg).id, ((x_3).ir_msg).type_, ((x_3).ir_msg).addr, (x_3).ir_msg_from, (x_3).ir_mshr_id, ((x_3).ir_by_victim).valid, ((x_3).ir_by_victim).data);
            countDone_fifoI2L_003 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoI2L_003 (Struct40 x_0);
        let x_1 = (full_fifoI2L_003);
        when (! (x_1), noAction);
        elt_fifoI2L_003 <= x_0;
        full_fifoI2L_003 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct40) deq_fifoI2L_003 ();
        let x_1 = (full_fifoI2L_003);
        when (x_1, noAction);
        let x_2 = (elt_fifoI2L_003);
        full_fifoI2L_003 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module93;
    method Action enq_fifoL2E_003 (Struct43 x_0);
    method ActionValue#(Struct43) deq_fifoL2E_003 ();
endinterface

module mkModule93
    (Module93);
    Reg#(Struct43) elt_fifoL2E_003 <- mkReg(unpack(0));
    Reg#(Bool) full_fifoL2E_003 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifoL2E_003 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifoL2E_003 <- mkReg(unpack(0));

    rule count_fifoL2E_003;

        let x_0 = (countDone_fifoL2E_003);
        when (! (x_0), noAction);
        let x_1 = (counter_fifoL2E_003);
        counter_fifoL2E_003 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifoL2E_003);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 =
            (elt_fifoL2E_003);
            $display ("-- LR fifoL2E_003: %b %x %b %x %x %x %b %x %x %b %x %b %x %b %x", ((x_3).lr_ir_pp).ir_is_rs_rel, (((x_3).lr_ir_pp).ir_msg).id, (((x_3).lr_ir_pp).ir_msg).type_, (((x_3).lr_ir_pp).ir_msg).addr, ((x_3).lr_ir_pp).ir_msg_from, ((x_3).lr_ir_pp).ir_mshr_id, (((x_3).lr_ir_pp).ir_by_victim).valid, (((x_3).lr_ir_pp).ir_by_victim).data, ((x_3).lr_ir).info_index, ((x_3).lr_ir).info_hit, ((x_3).lr_ir).info_way, ((x_3).lr_ir).edir_hit, ((x_3).lr_ir).edir_way, (((x_3).lr_ir).edir_slot).valid, (((x_3).lr_ir).edir_slot).data);
            countDone_fifoL2E_003 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifoL2E_003 (Struct43 x_0);
        let x_1 = (full_fifoL2E_003);
        when (! (x_1), noAction);
        elt_fifoL2E_003 <= x_0;
        full_fifoL2E_003 <= (Bool)'(True);
    endmethod

    method ActionValue#(Struct43) deq_fifoL2E_003 ();
        let x_1 = (full_fifoL2E_003);
        when (x_1, noAction);
        let x_2 = (elt_fifoL2E_003);
        full_fifoL2E_003 <= (Bool)'(False);
        return x_2;
    endmethod
endmodule

interface Module94;
    method Action enq_fifo0030 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0030 ();
endinterface

module mkModule94
    (Module94);
    Reg#(Vector#(2, Struct1)) elt_fifo0030 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0030 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0030 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0030 <- mkReg(True);
    Reg#(Bool) full_fifo0030 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0030 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0030 <- mkReg(unpack(0));

    rule count_fifo0030;

        let x_0 = (countDone_fifo0030);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0030);
        counter_fifo0030 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0030);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0030);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0030:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0030:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0030 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0030 (Struct1 x_0);
        let x_1 = (full_fifo0030);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0030);
        let x_3 = (enqP_fifo0030);
        let x_4 = (deqP_fifo0030);
        elt_fifo0030 <= update (x_2, x_3, x_0);
        empty_fifo0030 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0030 <= (x_4) == (x_5);
        enqP_fifo0030 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0030 ();
        let x_1 = (empty_fifo0030);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0030);
        let x_3 = (enqP_fifo0030);
        let x_4 = (deqP_fifo0030);
        full_fifo0030 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0030 <= (x_3) == (x_5);
        deqP_fifo0030 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module95;
    method Action enq_fifo0031 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0031 ();
endinterface

module mkModule95
    (Module95);
    Reg#(Vector#(2, Struct1)) elt_fifo0031 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0031 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0031 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0031 <- mkReg(True);
    Reg#(Bool) full_fifo0031 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0031 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0031 <- mkReg(unpack(0));

    rule count_fifo0031;

        let x_0 = (countDone_fifo0031);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0031);
        counter_fifo0031 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0031);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0031);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0031:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0031:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0031 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0031 (Struct1 x_0);
        let x_1 = (full_fifo0031);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0031);
        let x_3 = (enqP_fifo0031);
        let x_4 = (deqP_fifo0031);
        elt_fifo0031 <= update (x_2, x_3, x_0);
        empty_fifo0031 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0031 <= (x_4) == (x_5);
        enqP_fifo0031 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0031 ();
        let x_1 = (empty_fifo0031);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0031);
        let x_3 = (enqP_fifo0031);
        let x_4 = (deqP_fifo0031);
        full_fifo0031 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0031 <= (x_3) == (x_5);
        deqP_fifo0031 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module96;
    method Action enq_fifo0032 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0032 ();
endinterface

module mkModule96
    (Module96);
    Reg#(Vector#(2, Struct1)) elt_fifo0032 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo0032 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo0032 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo0032 <- mkReg(True);
    Reg#(Bool) full_fifo0032 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo0032 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo0032 <- mkReg(unpack(0));

    rule count_fifo0032;

        let x_0 = (countDone_fifo0032);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo0032);
        counter_fifo0032 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo0032);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo0032);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo0032:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo0032:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo0032 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo0032 (Struct1 x_0);
        let x_1 = (full_fifo0032);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0032);
        let x_3 = (enqP_fifo0032);
        let x_4 = (deqP_fifo0032);
        elt_fifo0032 <= update (x_2, x_3, x_0);
        empty_fifo0032 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo0032 <= (x_4) == (x_5);
        enqP_fifo0032 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo0032 ();
        let x_1 = (empty_fifo0032);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo0032);
        let x_3 = (enqP_fifo0032);
        let x_4 = (deqP_fifo0032);
        full_fifo0032 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo0032 <= (x_3) == (x_5);
        deqP_fifo0032 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module97;
    method Action enq_fifo00300 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00300 ();
endinterface

module mkModule97
    (Module97);
    Reg#(Vector#(2, Struct1)) elt_fifo00300 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00300 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00300 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00300 <- mkReg(True);
    Reg#(Bool) full_fifo00300 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00300 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00300 <- mkReg(unpack(0));

    rule count_fifo00300;

        let x_0 = (countDone_fifo00300);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00300);
        counter_fifo00300 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00300);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00300);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00300:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00300:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00300 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00300 (Struct1 x_0);
        let x_1 = (full_fifo00300);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00300);
        let x_3 = (enqP_fifo00300);
        let x_4 = (deqP_fifo00300);
        elt_fifo00300 <= update (x_2, x_3, x_0);
        empty_fifo00300 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00300 <= (x_4) == (x_5);
        enqP_fifo00300 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00300 ();
        let x_1 = (empty_fifo00300);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00300);
        let x_3 = (enqP_fifo00300);
        let x_4 = (deqP_fifo00300);
        full_fifo00300 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00300 <= (x_3) == (x_5);
        deqP_fifo00300 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module98;
    method Action enq_fifo00302 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00302 ();
endinterface

module mkModule98
    (Module98);
    Reg#(Vector#(2, Struct1)) elt_fifo00302 <- mkReg(unpack(0));
    Reg#(Bit#(1)) enqP_fifo00302 <- mkReg(unpack(0));
    Reg#(Bit#(1)) deqP_fifo00302 <- mkReg(unpack(0));
    Reg#(Bool) empty_fifo00302 <- mkReg(True);
    Reg#(Bool) full_fifo00302 <- mkReg(unpack(0));
    Reg#(Bool) countDone_fifo00302 <- mkReg(unpack(0));
    Reg#(Bit#(18)) counter_fifo00302 <- mkReg(unpack(0));

    rule count_fifo00302;

        let x_0 = (countDone_fifo00302);
        when (! (x_0), noAction);
        let x_1 = (counter_fifo00302);
        counter_fifo00302 <= (x_1) + ((Bit#(18))'(18'h1));
        let x_2 =
        (full_fifo00302);
        if (((x_1) == ((Bit#(18))'(18'h3ffff))) && (x_2)) begin
            let x_3 = (elt_fifo00302);
            Struct1 x_4 =
            ((x_3)[(Bit#(1))'(1'h1)]);
            $display ("-- MSG fifo00302:1 %x %b %x", (x_4).id, (x_4).type_, (x_4).addr);
            Struct1 x_5 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            $display ("-- MSG fifo00302:0 %x %b %x", (x_5).id, (x_5).type_, (x_5).addr);
            countDone_fifo00302 <= (Bool)'(True);
        end else begin

        end
    endrule

    method Action enq_fifo00302 (Struct1 x_0);
        let x_1 = (full_fifo00302);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00302);
        let x_3 = (enqP_fifo00302);
        let x_4 = (deqP_fifo00302);
        elt_fifo00302 <= update (x_2, x_3, x_0);
        empty_fifo00302 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_3) + ((Bit#(1))'(1'h1)));
        full_fifo00302 <= (x_4) == (x_5);
        enqP_fifo00302 <= x_5;
    endmethod

    method ActionValue#(Struct1) deq_fifo00302 ();
        let x_1 = (empty_fifo00302);
        when (! (x_1), noAction);
        let x_2 = (elt_fifo00302);
        let x_3 = (enqP_fifo00302);
        let x_4 = (deqP_fifo00302);
        full_fifo00302 <= (Bool)'(False);
        Bit#(1) x_5 = ((x_4) + ((Bit#(1))'(1'h1)));
        empty_fifo00302 <= (x_3) == (x_5);
        deqP_fifo00302 <= x_5;
        return (x_2)[x_4];
    endmethod
endmodule

interface Module99;
    method ActionValue#(Struct39) victims__003__findVictim (Bit#(64) x_0);
    method ActionValue#(Struct44) victims__003__getVictim (Bit#(2) x_0);
    method Action victims__003__setVictim (Struct48 x_0);
    method Action victims__003__registerVictim (Struct44 x_0);
    method ActionValue#(Struct44) victims__003__getFirstVictim ();
    method ActionValue#(Bool) victims__003__hasVictim ();
    method Action victims__003__setVictimRq (Struct49 x_0);
    method ActionValue#(Bit#(3)) victims__003__releaseVictim (Bit#(64) x_0);
endinterface

module mkModule99
    (Module99);
    Reg#(Vector#(4, Struct44)) victimRegs__003 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct39) victims__003__findVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__003);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_9 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            x_9 = Struct39 {valid : (Bool)'(True), data : (Bit#(2))'(2'h0)};
        end else begin
            Struct44 x_3 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_8 = ?;
            if (((x_3).victim_valid) && (((x_3).victim_addr) == (x_0)))
                begin
                x_8 = Struct39 {valid : (Bool)'(True), data :
                (Bit#(2))'(2'h1)};
            end else begin
                Struct44 x_4 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_7 = ?;
                if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                    begin
                    x_7 = Struct39 {valid : (Bool)'(True), data :
                    (Bit#(2))'(2'h2)};
                end else begin
                    Struct44 x_5 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_6 = ?;
                    if (((x_5).victim_valid) && (((x_5).victim_addr) ==
                        (x_0))) begin
                        x_6 = Struct39 {valid : (Bool)'(True), data :
                        (Bit#(2))'(2'h3)};
                    end else begin
                        x_6 = Struct39 {valid : (Bool)'(False), data :
                        unpack(0)};
                    end
                    x_7 = x_6;
                end
                x_8 = x_7;
            end
            x_9 = x_8;
        end
        return x_9;
    endmethod

    method ActionValue#(Struct44) victims__003__getVictim (Bit#(2) x_0);
        let x_1 = (victimRegs__003);
        return (x_1)[x_0];
    endmethod

    method Action victims__003__setVictim (Struct48 x_0);
        let x_1 = (victimRegs__003);
        Struct44 x_2 = ((x_1)[(x_0).victim_idx]);
        Struct44 x_3 = (Struct44 {victim_valid : (Bool)'(True), victim_addr :
        (x_2).victim_addr, victim_info : (x_0).victim_info, victim_value :
        (x_0).victim_value, victim_req : (x_2).victim_req});
        victimRegs__003 <= update (x_1, (x_0).victim_idx, x_3);
    endmethod

    method Action victims__003__registerVictim (Struct44 x_0);
        let x_1 = (victimRegs__003);
        Struct39 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_valid ? (Struct39 {valid :
        (Bool)'(False), data : unpack(0)}) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h0)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h1)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h2)}))) : (Struct39 {valid :
        (Bool)'(True), data : (Bit#(2))'(2'h3)})));
        when ((x_2).valid, noAction);
        Bit#(2) x_3 = ((x_2).data);
        victimRegs__003 <= update (x_1, x_3, x_0);
    endmethod

    method ActionValue#(Struct44) victims__003__getFirstVictim ();
        let x_1 = (victimRegs__003);
        Struct55 x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? (Struct55 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) : (Struct55 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method ActionValue#(Bool) victims__003__hasVictim ();
        let x_1 = (victimRegs__003);
        Bool x_2 = (((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h3)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_req).valid)) ? ((Bool)'(True)) :
        (((((x_1)[(Bit#(2))'(2'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(2))'(2'h0)]).victim_req).valid)) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        return x_2;
    endmethod

    method Action victims__003__setVictimRq (Struct49 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victimRegs__003);
        Struct44 x_4 =
        ((x_3)[(Bit#(2))'(2'h3)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct44 x_5 = (Struct44 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct5 {valid :
            (Bool)'(True), data : x_2}});
            victimRegs__003 <= update (x_3, (Bit#(2))'(2'h3), x_5);
        end else begin
            Struct44 x_6 =
            ((x_3)[(Bit#(2))'(2'h2)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct44 x_7 = (Struct44 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct5 {valid : (Bool)'(True), data :
                x_2}});
                victimRegs__003 <= update (x_3, (Bit#(2))'(2'h2), x_7);
            end else begin
                Struct44 x_8 =
                ((x_3)[(Bit#(2))'(2'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct44 x_9 = (Struct44 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct5 {valid :
                    (Bool)'(True), data : x_2}});
                    victimRegs__003 <= update (x_3, (Bit#(2))'(2'h1), x_9);
                end else begin
                    Struct44 x_10 =
                    ((x_3)[(Bit#(2))'(2'h0)]);
                    if (((x_10).victim_valid) && (((x_10).victim_addr) ==
                        (x_1))) begin
                        Struct44 x_11 = (Struct44 {victim_valid :
                        (x_10).victim_valid, victim_addr :
                        (x_10).victim_addr, victim_info : (x_10).victim_info,
                        victim_value : (x_10).victim_value, victim_req :
                        Struct5 {valid : (Bool)'(True), data :
                        x_2}});
                        victimRegs__003 <= update (x_3, (Bit#(2))'(2'h0),
                        x_11);
                    end else begin

                    end
                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) victims__003__releaseVictim (Bit#(64) x_0);
        let x_1 = (victimRegs__003);
        Struct44 x_2 =
        ((x_1)[(Bit#(2))'(2'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victimRegs__003 <= update (x_1, (Bit#(2))'(2'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct44 x_4 =
            ((x_1)[(Bit#(2))'(2'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victimRegs__003 <= update (x_1, (Bit#(2))'(2'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct44 x_6 =
                ((x_1)[(Bit#(2))'(2'h2)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victimRegs__003 <= update (x_1, (Bit#(2))'(2'h2),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct44 x_8 =
                    ((x_1)[(Bit#(2))'(2'h3)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victimRegs__003 <= update (x_1, (Bit#(2))'(2'h3),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod
endmodule

interface Module100;
    method Action rdReq_infoRam__003__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__003__3 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__003__3 ();
endinterface

module mkModule100 (Module100);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h7, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__003__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__003__3 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__003__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module101;
    method Action rdReq_infoRam__003__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__003__2 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__003__2 ();
endinterface

module mkModule101 (Module101);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h6, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__003__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__003__2 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__003__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module102;
    method Action rdReq_infoRam__003__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__003__1 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__003__1 ();
endinterface

module mkModule102 (Module102);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h5, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__003__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__003__1 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__003__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module103;
    method Action rdReq_infoRam__003__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__003__0 (Struct52 x_0);
    method ActionValue#(Struct50) rdResp_infoRam__003__0 ();
endinterface

module mkModule103 (Module103);
    RWBramCore#(Bit#(8), Struct50) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct50 {tag: 51'h4, value: Struct10 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 4'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__003__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__003__0 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct50) rdResp_infoRam__003__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module104;
    method Action rdReq_dataRam__003 (Bit#(10) x_0);
    method Action wrReq_dataRam__003 (Struct54 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__003 ();
endinterface

module mkModule104 (Module104);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__003 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__003 (Struct54 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__003 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module105;
    method Action rdReq_repRam__003 (Bit#(8) x_0);
    method Action wrReq_repRam__003 (Struct56 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__003 ();
endinterface

module mkModule105 (Module105);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h1, 8'h1, 8'h1, 8'h1);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__003 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__003 (Struct56 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__003 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module106;
    method ActionValue#(Struct45) getMSHR_003 (Bit#(3) x_0);
    method ActionValue#(Struct38) getPRqSlot_003 (Struct37 x_0);
    method ActionValue#(Struct38) getCRqSlot_003 (Struct37 x_0);
    method ActionValue#(Struct37) getWait_003 ();
    method Action registerUL_003 (Struct47 x_0);
    method Action registerDL_003 (Struct57 x_0);
    method Action canImm_003 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) setULImm_003 (Struct1 x_0);
    method Action transferUpDown_003 (Struct58 x_0);
    method Action addRs_003 (Struct7 x_0);
    method ActionValue#(Bit#(3)) getULReady_003 (Bit#(64) x_0);
    method ActionValue#(Struct59) getDLReady_003 ();
    method Action startRelease_003 (Bit#(3) x_0);
    method Action releaseMSHR_003 (Bit#(3) x_0);
endinterface

module mkModule106
    (Module106);
    Reg#(Vector#(6, Struct45)) rqs_003 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct45) getMSHR_003 (Bit#(3) x_0);
        let x_1 = (rqs_003);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct38) getPRqSlot_003 (Struct37 x_0);
        let x_1 = (rqs_003);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && (((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        || (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ?
        ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_8 = ((x_7).valid);
        Struct38 x_9 = (Struct38 {s_has_slot : (x_3) && (! (x_6)), s_conflict
        : x_8, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_10 = (update (x_1, x_4, Struct45 {m_status
            : (x_8 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_14 = ?;
            if (x_8) begin
                Bit#(3) x_11 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
                ((Bit#(3))'(3'h0)))) && (!
                ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h0)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h1)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h2)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h3)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h4)) : ((((!
                ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0))))
                && (! ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
                (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ?
                ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
                Struct45 x_12 = ((x_1)[x_11]);
                Vector#(6, Struct45) x_13 = (update (x_10, x_11, Struct45
                {m_status : (x_12).m_status, m_next : (x_8 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_12).m_next)), m_is_ul :
                (x_12).m_is_ul, m_msg : (x_12).m_msg, m_qidx : (x_12).m_qidx,
                m_rsb : (x_12).m_rsb, m_dl_rss_from : (x_12).m_dl_rss_from,
                m_dl_rss_recv : (x_12).m_dl_rss_recv, m_dl_rss :
                (x_12).m_dl_rss}));
                x_14 = x_13;
            end else begin
                x_14 = x_10;
            end
            rqs_003 <= x_14;
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct38) getCRqSlot_003 (Struct37 x_0);
        let x_1 = (rqs_003);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        Struct5 x_7 = (((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        Struct5 x_8 = (((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_9 = ((x_7).valid);
        Bool x_10 = ((x_8).valid);
        Bool x_11 = ((x_9) || (x_10));
        Struct38 x_12 = (Struct38 {s_has_slot : (x_3) && (! (x_6)),
        s_conflict : x_11, s_id :
        x_4});
        if ((x_3) && (! (x_6))) begin
            Vector#(6, Struct45) x_13 = (update (x_1, x_4, Struct45 {m_status
            : (x_11 ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h4))), m_next :
            Struct5 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul :
            unpack(0), m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb
            : unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv :
            unpack(0), m_dl_rss :
            unpack(0)}));
            let x_17 = ?;
            if (x_11) begin
                Bit#(3) x_14 = ((x_9 ? ((x_7).data) : ((x_8).data)));
                Struct45 x_15 = ((x_1)[x_14]);
                Vector#(6, Struct45) x_16 = (update (x_13, x_14, Struct45
                {m_status : (x_15).m_status, m_next : (x_11 ? (Struct5 {valid
                : (Bool)'(True), data : x_4}) : ((x_15).m_next)), m_is_ul :
                (x_15).m_is_ul, m_msg : (x_15).m_msg, m_qidx : (x_15).m_qidx,
                m_rsb : (x_15).m_rsb, m_dl_rss_from : (x_15).m_dl_rss_from,
                m_dl_rss_recv : (x_15).m_dl_rss_recv, m_dl_rss :
                (x_15).m_dl_rss}));
                x_17 = x_16;
            end else begin
                x_17 = x_13;
            end
            rqs_003 <= x_17;
        end else begin

        end
        return x_12;
    endmethod

    method ActionValue#(Struct37) getWait_003 ();
        let x_1 = (rqs_003);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h2)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h2)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((((! ((((x_1)[(Bit#(3))'(3'h4)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) ==
        (x_5))) || ((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5])))) ? ((Bool)'(True)) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) ||
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5]))))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        rqs_003 <= update (x_1, x_3, Struct45 {m_status : (Bit#(3))'(3'h4),
        m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg,
        m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : (x_4).m_dl_rss_recv, m_dl_rss :
        (x_4).m_dl_rss});
        Struct37 x_7 = (Struct37 {r_id : x_3, r_msg : (x_4).m_msg, r_msg_from
        : (x_4).m_qidx});
        return x_7;
    endmethod

    method Action registerUL_003 (Struct47 x_0);
        let x_1 = (rqs_003);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_003 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_003 (Struct57 x_0);
        let x_1 = (rqs_003);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_003 <= update (x_1, x_2, x_4);
    endmethod

    method Action canImm_003 (Bit#(64) x_0);
        let x_1 = (rqs_003);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
    endmethod

    method ActionValue#(Bit#(3)) setULImm_003 (Struct1 x_0);
        let x_1 = (rqs_003);
        Struct5 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(3))'(3'h0)) ? (Struct5 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct5 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Bit#(64) x_4 = ((x_0).addr);
        Struct5 x_5 = (((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h0)))) && (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) ==
        (x_4)) ? (Struct5 {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((! ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : (((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h0)))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_4)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_5).valid), noAction);
        Vector#(6, Struct45) x_6 = (update (x_1, x_3, Struct45 {m_status :
        (Bit#(3))'(3'h5), m_next : Struct5 {valid : (Bool)'(False), data :
        unpack(0)}, m_is_ul : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)}));
        rqs_003 <= x_6;
        return x_3;
    endmethod

    method Action transferUpDown_003 (Struct58 x_0);
        let x_1 = (rqs_003);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct45 x_3 = ((x_1)[x_2]);
        Struct45 x_4 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_003 <= update (x_1, x_2, x_4);
    endmethod

    method Action addRs_003 (Struct7 x_0);
        let x_1 = (rqs_003);
        Bit#(64) x_2 = (((x_0).r_msg).addr);
        Struct5 x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_3).valid, noAction);
        Bit#(3) x_4 = ((x_3).data);
        Struct45 x_5 = ((x_1)[x_4]);
        Struct45 x_6 = (Struct45 {m_status : (x_5).m_status, m_next :
        (x_5).m_next, m_is_ul : (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx :
        (x_5).m_qidx, m_rsb : (x_5).m_rsb, m_dl_rss_from :
        (x_5).m_dl_rss_from, m_dl_rss_recv : ((x_5).m_dl_rss_recv) |
        (((Bit#(4))'(4'h1)) << ((x_0).r_midx)), m_dl_rss : update
        ((x_5).m_dl_rss, (x_0).r_midx, (x_0).r_msg)});
        rqs_003 <= update (x_1, x_4, x_6);
    endmethod

    method ActionValue#(Bit#(3)) getULReady_003 (Bit#(64) x_0);
        let x_1 = (rqs_003);
        Bool x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_0))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_0)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_0)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_2), noAction);
        Struct5 x_3 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) <
        ((Bit#(3))'(3'h4)))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) < ((Bit#(3))'(3'h4)))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when (! ((x_3).valid), noAction);
        Struct5 x_4 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) &&
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))));
        when ((x_4).valid, noAction);
        Bit#(3) x_5 = ((x_4).data);
        return x_5;
    endmethod

    method ActionValue#(Struct59) getDLReady_003 ();
        let x_1 = (rqs_003);
        Struct5 x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h5))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h0)}) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h1)}) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h2)}) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h3)}) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h4)}) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h5))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? (Struct5 {valid :
        (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        Struct45 x_4 = ((x_1)[x_3]);
        Bit#(64) x_5 = (((x_4).m_msg).addr);
        Bool x_6 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h4))) || ((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(3))'(3'h6)))) && ((! (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)
        == (x_5))) && ((((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr)[12:5]) ==
        ((x_5)[12:5]))) ? ((Bool)'(True)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h4))) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(3))'(3'h6)))) && ((!
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5))) &&
        ((((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr)[12:5]) == ((x_5)[12:5])))
        ? ((Bool)'(True)) : ((Bool)'(False))))))))))))));
        when (! (x_6), noAction);
        Struct59 x_7 = (Struct59 {r_id : x_3, r_addr : x_5});
        return x_7;
    endmethod

    method Action startRelease_003 (Bit#(3) x_0);
        let x_1 = (rqs_003);
        Struct45 x_2 = ((x_1)[x_0]);
        Struct45 x_3 = (Struct45 {m_status : (Bit#(3))'(3'h6), m_next :
        (x_2).m_next, m_is_ul : (x_2).m_is_ul, m_msg : (x_2).m_msg, m_qidx :
        (x_2).m_qidx, m_rsb : (x_2).m_rsb, m_dl_rss_from :
        (x_2).m_dl_rss_from, m_dl_rss_recv : (x_2).m_dl_rss_recv, m_dl_rss :
        (x_2).m_dl_rss});
        rqs_003 <= update (x_1, x_0, x_3);
    endmethod

    method Action releaseMSHR_003 (Bit#(3) x_0);
        let x_1 = (rqs_003);
        Struct45 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct45) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct45 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct45) x_6 = (update (x_3, x_4, Struct45 {m_status
            : (Bit#(3))'(3'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_003 <= x_7;
    endmethod
endmodule

interface Module107;

endinterface

module mkModule107#(function ActionValue#(Struct1) deq_fifo0030(),
    function ActionValue#(Struct1) deq_fifo0020(),
    function ActionValue#(Struct1) deq_fifo0010(),
    function Action enq_fifoCRqInput_00(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0000())
    (Module107);
    Reg#(Bit#(2)) rr_cRq4_00 <- mkReg(unpack(0));

    rule inc_rr_cRq4_00;

        let x_0 = (rr_cRq4_00);
        rr_cRq4_00 <= (x_0) + ((Bit#(2))'(2'h1));
    endrule

    rule accept0_cRq4_00;
        $display ("Rule fired: accept0_cRq4_00 at %t", $time);
        let x_0 = (rr_cRq4_00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 <- deq_fifo0000();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h0))}});
        let x_3 <- enq_fifoCRqInput_00(x_2);
    endrule

    rule accept1_cRq4_00;
        $display ("Rule fired: accept1_cRq4_00 at %t", $time);
        let x_0 = (rr_cRq4_00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 <- deq_fifo0010();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h1))}});
        let x_3 <- enq_fifoCRqInput_00(x_2);
    endrule

    rule accept2_cRq4_00;
        $display ("Rule fired: accept2_cRq4_00 at %t", $time);
        let x_0 = (rr_cRq4_00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 <- deq_fifo0020();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h2))}});
        let x_3 <- enq_fifoCRqInput_00(x_2);
    endrule

    rule accept3_cRq4_00;
        $display ("Rule fired: accept3_cRq4_00 at %t", $time);
        let x_0 = (rr_cRq4_00);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 <- deq_fifo0030();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h3))}});
        let x_3 <- enq_fifoCRqInput_00(x_2);
    endrule

    // No methods in this module
endmodule

interface Module108;

endinterface

module mkModule108#(function ActionValue#(Struct1) deq_fifo0031(),
    function ActionValue#(Struct1) deq_fifo0021(),
    function ActionValue#(Struct1) deq_fifo0011(),
    function Action enq_fifoCRsInput_00(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0001())
    (Module108);
    Reg#(Bit#(2)) rr_cRs4_00 <- mkReg(unpack(0));

    rule inc_rr_cRs4_00;

        let x_0 = (rr_cRs4_00);
        rr_cRs4_00 <= (x_0) + ((Bit#(2))'(2'h1));
    endrule

    rule accept0_cRs4_00;
        $display ("Rule fired: accept0_cRs4_00 at %t", $time);
        let x_0 = (rr_cRs4_00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 <- deq_fifo0001();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h1)),((Bit#(2))'(2'h0))}});
        let x_3 <- enq_fifoCRsInput_00(x_2);
    endrule

    rule accept1_cRs4_00;
        $display ("Rule fired: accept1_cRs4_00 at %t", $time);
        let x_0 = (rr_cRs4_00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 <- deq_fifo0011();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h1)),((Bit#(2))'(2'h1))}});
        let x_3 <- enq_fifoCRsInput_00(x_2);
    endrule

    rule accept2_cRs4_00;
        $display ("Rule fired: accept2_cRs4_00 at %t", $time);
        let x_0 = (rr_cRs4_00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 <- deq_fifo0021();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h1)),((Bit#(2))'(2'h2))}});
        let x_3 <- enq_fifoCRsInput_00(x_2);
    endrule

    rule accept3_cRs4_00;
        $display ("Rule fired: accept3_cRs4_00 at %t", $time);
        let x_0 = (rr_cRs4_00);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 <- deq_fifo0031();
        Struct2 x_2 = (Struct2 {in_msg : x_1, in_msg_from :
        {((Bit#(2))'(2'h1)),((Bit#(2))'(2'h3))}});
        let x_3 <- enq_fifoCRsInput_00(x_2);
    endrule

    // No methods in this module
endmodule

interface Module109;

endinterface

module mkModule109#(function Action enq_fifoPInput_00(Struct2 _),
    function ActionValue#(Struct1) deq_fifo002())
    (Module109);

    rule parent_convert_00;
        $display ("Rule fired: parent_convert_00 at %t", $time);
        let x_0 <- deq_fifo002();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}});
        let x_2 <- enq_fifoPInput_00(x_1);
    endrule

    // No methods in this module
endmodule

interface Module110;
    method Action makeEnq_parentChildren00 (Struct19 x_0);
    method Action broadcast_parentChildren00 (Struct22 x_0);
endinterface

module mkModule110#(function Action enq_fifo0002(Struct1 _),
    function Action enq_fifo0012(Struct1 _),
    function Action enq_fifo0022(Struct1 _),
    function Action enq_fifo0032(Struct1 _),
    function Action enq_fifo001(Struct1 _),
    function Action enq_fifo000(Struct1 _))
    (Module110);

    // No rules in this module

    method Action makeEnq_parentChildren00 (Struct19 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo000((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo001((x_0).enq_msg);
            end else begin
                Bit#(2) x_3 = ((x_0).enq_ch_idx);
                Struct1 x_4 =
                ((x_0).enq_msg);
                if ((x_3) == ((Bit#(2))'(2'h3))) begin
                    let x_5 <- enq_fifo0032(x_4);
                end else
                    begin
                    if ((x_3) == ((Bit#(2))'(2'h2))) begin
                        let x_6 <- enq_fifo0022(x_4);
                    end else
                        begin
                        if ((x_3) == ((Bit#(2))'(2'h1))) begin
                            let x_7 <- enq_fifo0012(x_4);
                        end else
                            begin
                            if ((x_3) == ((Bit#(2))'(2'h0))) begin
                                let x_8 <- enq_fifo0002(x_4);
                            end else begin

                            end
                        end
                    end
                end
            end
        end
    endmethod

    method Action broadcast_parentChildren00 (Struct22 x_0);
        Bit#(4) x_1 = ((x_0).cs_inds);
        Struct1 x_2 =
        ((x_0).cs_msg);
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == (x_1))
            begin
            let x_3 <- enq_fifo0032(x_2);
        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == (x_1))
            begin
            let x_5 <- enq_fifo0022(x_2);
        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == (x_1))
            begin
            let x_7 <- enq_fifo0012(x_2);
        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == (x_1))
            begin
            let x_9 <- enq_fifo0002(x_2);
        end else begin

        end
    endmethod
endmodule

interface Module111;
    method Action repGetRq__00 (Bit#(9) x_0);
    method ActionValue#(Vector#(16, Bit#(8))) repGetRs__00 ();
    method Action repAccess__00 (Struct32 x_0);
endinterface

module mkModule111#(function Action wrReq_repRam__00(Struct36 _),
    function ActionValue#(Vector#(16, Bit#(8))) rdResp_repRam__00(),
    function Action rdReq_repRam__00(Bit#(9) _))
    (Module111);

    // No rules in this module

    method Action repGetRq__00 (Bit#(9) x_0);
        let x_1 <- rdReq_repRam__00(x_0);
    endmethod

    method ActionValue#(Vector#(16, Bit#(8))) repGetRs__00 ();
        let x_1 <- rdResp_repRam__00();
        return x_1;
    endmethod

    method Action repAccess__00 (Struct32 x_0);
        Vector#(16, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(4))'(4'hf)]) +
        (((((x_1)[(Bit#(4))'(4'hf)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(4))'(4'hf)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_3 = (update (x_1, (Bit#(4))'(4'hf),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(4))'(4'he)]) +
        (((((x_3)[(Bit#(4))'(4'he)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(4))'(4'he)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_5 = (update (x_3, (Bit#(4))'(4'he),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(4))'(4'hd)]) +
        (((((x_5)[(Bit#(4))'(4'hd)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(4))'(4'hd)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_7 = (update (x_5, (Bit#(4))'(4'hd),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(4))'(4'hc)]) +
        (((((x_7)[(Bit#(4))'(4'hc)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(4))'(4'hc)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_9 = (update (x_7, (Bit#(4))'(4'hc),
        x_8));
        Bit#(8) x_10 = (((x_9)[(Bit#(4))'(4'hb)]) +
        (((((x_9)[(Bit#(4))'(4'hb)]) == ((Bit#(8))'(8'h0))) ||
        (((x_9)[(Bit#(4))'(4'hb)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_11 = (update (x_9, (Bit#(4))'(4'hb),
        x_10));
        Bit#(8) x_12 = (((x_11)[(Bit#(4))'(4'ha)]) +
        (((((x_11)[(Bit#(4))'(4'ha)]) == ((Bit#(8))'(8'h0))) ||
        (((x_11)[(Bit#(4))'(4'ha)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_13 = (update (x_11, (Bit#(4))'(4'ha),
        x_12));
        Bit#(8) x_14 = (((x_13)[(Bit#(4))'(4'h9)]) +
        (((((x_13)[(Bit#(4))'(4'h9)]) == ((Bit#(8))'(8'h0))) ||
        (((x_13)[(Bit#(4))'(4'h9)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_15 = (update (x_13, (Bit#(4))'(4'h9),
        x_14));
        Bit#(8) x_16 = (((x_15)[(Bit#(4))'(4'h8)]) +
        (((((x_15)[(Bit#(4))'(4'h8)]) == ((Bit#(8))'(8'h0))) ||
        (((x_15)[(Bit#(4))'(4'h8)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_17 = (update (x_15, (Bit#(4))'(4'h8),
        x_16));
        Bit#(8) x_18 = (((x_17)[(Bit#(4))'(4'h7)]) +
        (((((x_17)[(Bit#(4))'(4'h7)]) == ((Bit#(8))'(8'h0))) ||
        (((x_17)[(Bit#(4))'(4'h7)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_19 = (update (x_17, (Bit#(4))'(4'h7),
        x_18));
        Bit#(8) x_20 = (((x_19)[(Bit#(4))'(4'h6)]) +
        (((((x_19)[(Bit#(4))'(4'h6)]) == ((Bit#(8))'(8'h0))) ||
        (((x_19)[(Bit#(4))'(4'h6)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_21 = (update (x_19, (Bit#(4))'(4'h6),
        x_20));
        Bit#(8) x_22 = (((x_21)[(Bit#(4))'(4'h5)]) +
        (((((x_21)[(Bit#(4))'(4'h5)]) == ((Bit#(8))'(8'h0))) ||
        (((x_21)[(Bit#(4))'(4'h5)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_23 = (update (x_21, (Bit#(4))'(4'h5),
        x_22));
        Bit#(8) x_24 = (((x_23)[(Bit#(4))'(4'h4)]) +
        (((((x_23)[(Bit#(4))'(4'h4)]) == ((Bit#(8))'(8'h0))) ||
        (((x_23)[(Bit#(4))'(4'h4)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_25 = (update (x_23, (Bit#(4))'(4'h4),
        x_24));
        Bit#(8) x_26 = (((x_25)[(Bit#(4))'(4'h3)]) +
        (((((x_25)[(Bit#(4))'(4'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_25)[(Bit#(4))'(4'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_27 = (update (x_25, (Bit#(4))'(4'h3),
        x_26));
        Bit#(8) x_28 = (((x_27)[(Bit#(4))'(4'h2)]) +
        (((((x_27)[(Bit#(4))'(4'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_27)[(Bit#(4))'(4'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_29 = (update (x_27, (Bit#(4))'(4'h2),
        x_28));
        Bit#(8) x_30 = (((x_29)[(Bit#(4))'(4'h1)]) +
        (((((x_29)[(Bit#(4))'(4'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_29)[(Bit#(4))'(4'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_31 = (update (x_29, (Bit#(4))'(4'h1),
        x_30));
        Bit#(8) x_32 = (((x_31)[(Bit#(4))'(4'h0)]) +
        (((((x_31)[(Bit#(4))'(4'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_31)[(Bit#(4))'(4'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_33 = (update (x_31, (Bit#(4))'(4'h0),
        x_32));
        let x_36 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(16, Bit#(8)) x_34 = (update (x_33, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_36 = x_34;
        end else begin
            Vector#(16, Bit#(8)) x_35 = (update (x_33, (x_0).acc_way,
            (Bit#(8))'(8'h0)));
            x_36 = x_35;
        end
        Struct36 x_37 = (Struct36 {addr : (x_0).acc_index, datain :
        x_36});
        let x_38 <- wrReq_repRam__00(x_37);
    endmethod
endmodule

interface Module112;

endinterface

module mkModule112#(function Action enq_fifoCRqInput_000(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00000())
    (Module112);

    rule child_convert_000;
        $display ("Rule fired: child_convert_000 at %t", $time);
        let x_0 <- deq_fifo00000();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h0))}});
        let x_2 <- enq_fifoCRqInput_000(x_1);
    endrule

    // No methods in this module
endmodule

interface Module113;

endinterface

module mkModule113#(function Action enq_fifoPInput_000(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0002())
    (Module113);

    rule parent_convert_000;
        $display ("Rule fired: parent_convert_000 at %t", $time);
        let x_0 <- deq_fifo0002();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}});
        let x_2 <- enq_fifoPInput_000(x_1);
    endrule

    // No methods in this module
endmodule

interface Module114;
    method Action makeEnq_parentChildren000 (Struct19 x_0);
endinterface

module mkModule114#(function Action enq_fifo00002(Struct1 _),
    function Action enq_fifo0001(Struct1 _),
    function Action enq_fifo0000(Struct1 _))
    (Module114);

    // No rules in this module

    method Action makeEnq_parentChildren000 (Struct19 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo0000((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo0001((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo00002(x_3);
            end
        end
    endmethod
endmodule

interface Module115;
    method Action repGetRq__000 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__000 ();
    method Action repAccess__000 (Struct53 x_0);
endinterface

module mkModule115#(function Action wrReq_repRam__000(Struct56 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__000(),
    function Action rdReq_repRam__000(Bit#(8) _))
    (Module115);

    // No rules in this module

    method Action repGetRq__000 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__000(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__000 ();
        let x_1 <- rdResp_repRam__000();
        return x_1;
    endmethod

    method Action repAccess__000 (Struct53 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h0)));
            x_12 = x_11;
        end
        Struct56 x_13 = (Struct56 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__000(x_13);
    endmethod
endmodule

interface Module116;

endinterface

module mkModule116#(function Action enq_fifoCRqInput_001(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00100())
    (Module116);

    rule child_convert_001;
        $display ("Rule fired: child_convert_001 at %t", $time);
        let x_0 <- deq_fifo00100();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h0))}});
        let x_2 <- enq_fifoCRqInput_001(x_1);
    endrule

    // No methods in this module
endmodule

interface Module117;

endinterface

module mkModule117#(function Action enq_fifoPInput_001(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0012())
    (Module117);

    rule parent_convert_001;
        $display ("Rule fired: parent_convert_001 at %t", $time);
        let x_0 <- deq_fifo0012();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h2)),((Bit#(2))'(2'h1))}});
        let x_2 <- enq_fifoPInput_001(x_1);
    endrule

    // No methods in this module
endmodule

interface Module118;
    method Action makeEnq_parentChildren001 (Struct19 x_0);
endinterface

module mkModule118#(function Action enq_fifo00102(Struct1 _),
    function Action enq_fifo0011(Struct1 _),
    function Action enq_fifo0010(Struct1 _))
    (Module118);

    // No rules in this module

    method Action makeEnq_parentChildren001 (Struct19 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo0010((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo0011((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo00102(x_3);
            end
        end
    endmethod
endmodule

interface Module119;
    method Action repGetRq__001 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__001 ();
    method Action repAccess__001 (Struct53 x_0);
endinterface

module mkModule119#(function Action wrReq_repRam__001(Struct56 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__001(),
    function Action rdReq_repRam__001(Bit#(8) _))
    (Module119);

    // No rules in this module

    method Action repGetRq__001 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__001(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__001 ();
        let x_1 <- rdResp_repRam__001();
        return x_1;
    endmethod

    method Action repAccess__001 (Struct53 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h0)));
            x_12 = x_11;
        end
        Struct56 x_13 = (Struct56 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__001(x_13);
    endmethod
endmodule

interface Module120;

endinterface

module mkModule120#(function Action enq_fifoCRqInput_002(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00200())
    (Module120);

    rule child_convert_002;
        $display ("Rule fired: child_convert_002 at %t", $time);
        let x_0 <- deq_fifo00200();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h0))}});
        let x_2 <- enq_fifoCRqInput_002(x_1);
    endrule

    // No methods in this module
endmodule

interface Module121;

endinterface

module mkModule121#(function Action enq_fifoPInput_002(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0022())
    (Module121);

    rule parent_convert_002;
        $display ("Rule fired: parent_convert_002 at %t", $time);
        let x_0 <- deq_fifo0022();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h2)),((Bit#(2))'(2'h2))}});
        let x_2 <- enq_fifoPInput_002(x_1);
    endrule

    // No methods in this module
endmodule

interface Module122;
    method Action makeEnq_parentChildren002 (Struct19 x_0);
endinterface

module mkModule122#(function Action enq_fifo00202(Struct1 _),
    function Action enq_fifo0021(Struct1 _),
    function Action enq_fifo0020(Struct1 _))
    (Module122);

    // No rules in this module

    method Action makeEnq_parentChildren002 (Struct19 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo0020((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo0021((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo00202(x_3);
            end
        end
    endmethod
endmodule

interface Module123;
    method Action repGetRq__002 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__002 ();
    method Action repAccess__002 (Struct53 x_0);
endinterface

module mkModule123#(function Action wrReq_repRam__002(Struct56 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__002(),
    function Action rdReq_repRam__002(Bit#(8) _))
    (Module123);

    // No rules in this module

    method Action repGetRq__002 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__002(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__002 ();
        let x_1 <- rdResp_repRam__002();
        return x_1;
    endmethod

    method Action repAccess__002 (Struct53 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h0)));
            x_12 = x_11;
        end
        Struct56 x_13 = (Struct56 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__002(x_13);
    endmethod
endmodule

interface Module124;

endinterface

module mkModule124#(function Action enq_fifoCRqInput_003(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00300())
    (Module124);

    rule child_convert_003;
        $display ("Rule fired: child_convert_003 at %t", $time);
        let x_0 <- deq_fifo00300();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h0)),((Bit#(2))'(2'h0))}});
        let x_2 <- enq_fifoCRqInput_003(x_1);
    endrule

    // No methods in this module
endmodule

interface Module125;

endinterface

module mkModule125#(function Action enq_fifoPInput_003(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0032())
    (Module125);

    rule parent_convert_003;
        $display ("Rule fired: parent_convert_003 at %t", $time);
        let x_0 <- deq_fifo0032();
        Struct2 x_1 = (Struct2 {in_msg : x_0, in_msg_from :
        {((Bit#(2))'(2'h2)),((Bit#(2))'(2'h3))}});
        let x_2 <- enq_fifoPInput_003(x_1);
    endrule

    // No methods in this module
endmodule

interface Module126;
    method Action makeEnq_parentChildren003 (Struct19 x_0);
endinterface

module mkModule126#(function Action enq_fifo00302(Struct1 _),
    function Action enq_fifo0031(Struct1 _),
    function Action enq_fifo0030(Struct1 _))
    (Module126);

    // No rules in this module

    method Action makeEnq_parentChildren003 (Struct19 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo0030((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo0031((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo00302(x_3);
            end
        end
    endmethod
endmodule

interface Module127;
    method Action repGetRq__003 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__003 ();
    method Action repAccess__003 (Struct53 x_0);
endinterface

module mkModule127#(function Action wrReq_repRam__003(Struct56 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__003(),
    function Action rdReq_repRam__003(Bit#(8) _))
    (Module127);

    // No rules in this module

    method Action repGetRq__003 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__003(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__003 ();
        let x_1 <- rdResp_repRam__003();
        return x_1;
    endmethod

    method Action repAccess__003 (Struct53 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h0)));
            x_12 = x_11;
        end
        Struct56 x_13 = (Struct56 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__003(x_13);
    endmethod
endmodule

interface Module128;
    method Action cache__00__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct9) cache__00__infoRsValueRq (Bit#(64) x_0);
    method ActionValue#(Vector#(4, Bit#(64))) cache__00__valueRsLineRq
    (Struct17 x_0);
endinterface

module mkModule128#(function Action wrReq_dataRam__00(Struct34 _),
    function Action wrReq_edirRam__00__7(Struct33 _),
    function Action wrReq_edirRam__00__6(Struct33 _),
    function Action wrReq_edirRam__00__5(Struct33 _),
    function Action wrReq_edirRam__00__4(Struct33 _),
    function Action wrReq_edirRam__00__3(Struct33 _),
    function Action wrReq_edirRam__00__2(Struct33 _),
    function Action wrReq_edirRam__00__1(Struct33 _),
    function Action wrReq_edirRam__00__0(Struct33 _),
    function Action repAccess__00(Struct32 _),
    function Action victims__00__registerVictim(Struct13 _),
    function Action wrReq_infoRam__00__15(Struct31 _),
    function Action wrReq_infoRam__00__14(Struct31 _),
    function Action wrReq_infoRam__00__13(Struct31 _),
    function Action wrReq_infoRam__00__12(Struct31 _),
    function Action wrReq_infoRam__00__11(Struct31 _),
    function Action wrReq_infoRam__00__10(Struct31 _),
    function Action wrReq_infoRam__00__9(Struct31 _),
    function Action wrReq_infoRam__00__8(Struct31 _),
    function Action wrReq_infoRam__00__7(Struct31 _),
    function Action wrReq_infoRam__00__6(Struct31 _),
    function Action wrReq_infoRam__00__5(Struct31 _),
    function Action wrReq_infoRam__00__4(Struct31 _),
    function Action wrReq_infoRam__00__3(Struct31 _),
    function Action wrReq_infoRam__00__2(Struct31 _),
    function Action wrReq_infoRam__00__1(Struct31 _),
    function Action wrReq_infoRam__00__0(Struct31 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__00(),
    function Action rdReq_dataRam__00(Bit#(13) _),
    function ActionValue#(Vector#(16, Bit#(8))) repGetRs__00(),
    function ActionValue#(Struct28) rdResp_edirRam__00__7(),
    function ActionValue#(Struct28) rdResp_edirRam__00__6(),
    function ActionValue#(Struct28) rdResp_edirRam__00__5(),
    function ActionValue#(Struct28) rdResp_edirRam__00__4(),
    function ActionValue#(Struct28) rdResp_edirRam__00__3(),
    function ActionValue#(Struct28) rdResp_edirRam__00__2(),
    function ActionValue#(Struct28) rdResp_edirRam__00__1(),
    function ActionValue#(Struct28) rdResp_edirRam__00__0(),
    function ActionValue#(Struct26) rdResp_infoRam__00__15(),
    function ActionValue#(Struct26) rdResp_infoRam__00__14(),
    function ActionValue#(Struct26) rdResp_infoRam__00__13(),
    function ActionValue#(Struct26) rdResp_infoRam__00__12(),
    function ActionValue#(Struct26) rdResp_infoRam__00__11(),
    function ActionValue#(Struct26) rdResp_infoRam__00__10(),
    function ActionValue#(Struct26) rdResp_infoRam__00__9(),
    function ActionValue#(Struct26) rdResp_infoRam__00__8(),
    function ActionValue#(Struct26) rdResp_infoRam__00__7(),
    function ActionValue#(Struct26) rdResp_infoRam__00__6(),
    function ActionValue#(Struct26) rdResp_infoRam__00__5(),
    function ActionValue#(Struct26) rdResp_infoRam__00__4(),
    function ActionValue#(Struct26) rdResp_infoRam__00__3(),
    function ActionValue#(Struct26) rdResp_infoRam__00__2(),
    function ActionValue#(Struct26) rdResp_infoRam__00__1(),
    function ActionValue#(Struct26) rdResp_infoRam__00__0(),
    function Action repGetRq__00(Bit#(9) _),
    function Action rdReq_edirRam__00__7(Bit#(9) _),
    function Action rdReq_edirRam__00__6(Bit#(9) _),
    function Action rdReq_edirRam__00__5(Bit#(9) _),
    function Action rdReq_edirRam__00__4(Bit#(9) _),
    function Action rdReq_edirRam__00__3(Bit#(9) _),
    function Action rdReq_edirRam__00__2(Bit#(9) _),
    function Action rdReq_edirRam__00__1(Bit#(9) _),
    function Action rdReq_edirRam__00__0(Bit#(9) _),
    function Action rdReq_infoRam__00__15(Bit#(9) _),
    function Action rdReq_infoRam__00__14(Bit#(9) _),
    function Action rdReq_infoRam__00__13(Bit#(9) _),
    function Action rdReq_infoRam__00__12(Bit#(9) _),
    function Action rdReq_infoRam__00__11(Bit#(9) _),
    function Action rdReq_infoRam__00__10(Bit#(9) _),
    function Action rdReq_infoRam__00__9(Bit#(9) _),
    function Action rdReq_infoRam__00__8(Bit#(9) _),
    function Action rdReq_infoRam__00__7(Bit#(9) _),
    function Action rdReq_infoRam__00__6(Bit#(9) _),
    function Action rdReq_infoRam__00__5(Bit#(9) _),
    function Action rdReq_infoRam__00__4(Bit#(9) _),
    function Action rdReq_infoRam__00__3(Bit#(9) _),
    function Action rdReq_infoRam__00__2(Bit#(9) _),
    function Action rdReq_infoRam__00__1(Bit#(9) _),
    function Action rdReq_infoRam__00__0(Bit#(9) _))
    (Module128);

    // No rules in this module

    method Action cache__00__infoRq (Bit#(64) x_0);
        Bit#(9) x_1 = ((x_0)[13:5]);
        let x_2 <- rdReq_infoRam__00__0(x_1);
        let x_3 <- rdReq_infoRam__00__1(x_1);
        let x_4 <- rdReq_infoRam__00__2(x_1);
        let x_5 <- rdReq_infoRam__00__3(x_1);
        let x_6 <- rdReq_infoRam__00__4(x_1);
        let x_7 <- rdReq_infoRam__00__5(x_1);
        let x_8 <- rdReq_infoRam__00__6(x_1);
        let x_9 <- rdReq_infoRam__00__7(x_1);
        let x_10 <- rdReq_infoRam__00__8(x_1);
        let x_11 <- rdReq_infoRam__00__9(x_1);
        let x_12 <- rdReq_infoRam__00__10(x_1);
        let x_13 <- rdReq_infoRam__00__11(x_1);
        let x_14 <- rdReq_infoRam__00__12(x_1);
        let x_15 <- rdReq_infoRam__00__13(x_1);
        let x_16 <- rdReq_infoRam__00__14(x_1);
        let x_17 <- rdReq_infoRam__00__15(x_1);
        let x_18 <- rdReq_edirRam__00__0(x_1);
        let x_19 <- rdReq_edirRam__00__1(x_1);
        let x_20 <- rdReq_edirRam__00__2(x_1);
        let x_21 <- rdReq_edirRam__00__3(x_1);
        let x_22 <- rdReq_edirRam__00__4(x_1);
        let x_23 <- rdReq_edirRam__00__5(x_1);
        let x_24 <- rdReq_edirRam__00__6(x_1);
        let x_25 <- rdReq_edirRam__00__7(x_1);
        let x_26 <- repGetRq__00(x_1);
    endmethod

    method ActionValue#(Struct9) cache__00__infoRsValueRq (Bit#(64) x_0);
        Bit#(50) x_1 = ((x_0)[63:14]);
        Bit#(9) x_2 = ((x_0)[13:5]);
        Vector#(16, Struct26) x_3 = (unpack(0));
        let x_4 <- rdResp_infoRam__00__0();
        Vector#(16, Struct26) x_5 = (update (x_3, (Bit#(4))'(4'h0), x_4));
        let x_6 <- rdResp_infoRam__00__1();
        Vector#(16, Struct26) x_7 = (update (x_5, (Bit#(4))'(4'h1), x_6));
        let x_8 <- rdResp_infoRam__00__2();
        Vector#(16, Struct26) x_9 = (update (x_7, (Bit#(4))'(4'h2), x_8));
        let x_10 <- rdResp_infoRam__00__3();
        Vector#(16, Struct26) x_11 = (update (x_9, (Bit#(4))'(4'h3),
        x_10));
        let x_12 <- rdResp_infoRam__00__4();
        Vector#(16, Struct26) x_13 = (update (x_11, (Bit#(4))'(4'h4),
        x_12));
        let x_14 <- rdResp_infoRam__00__5();
        Vector#(16, Struct26) x_15 = (update (x_13, (Bit#(4))'(4'h5),
        x_14));
        let x_16 <- rdResp_infoRam__00__6();
        Vector#(16, Struct26) x_17 = (update (x_15, (Bit#(4))'(4'h6),
        x_16));
        let x_18 <- rdResp_infoRam__00__7();
        Vector#(16, Struct26) x_19 = (update (x_17, (Bit#(4))'(4'h7),
        x_18));
        let x_20 <- rdResp_infoRam__00__8();
        Vector#(16, Struct26) x_21 = (update (x_19, (Bit#(4))'(4'h8),
        x_20));
        let x_22 <- rdResp_infoRam__00__9();
        Vector#(16, Struct26) x_23 = (update (x_21, (Bit#(4))'(4'h9),
        x_22));
        let x_24 <- rdResp_infoRam__00__10();
        Vector#(16, Struct26) x_25 = (update (x_23, (Bit#(4))'(4'ha),
        x_24));
        let x_26 <- rdResp_infoRam__00__11();
        Vector#(16, Struct26) x_27 = (update (x_25, (Bit#(4))'(4'hb),
        x_26));
        let x_28 <- rdResp_infoRam__00__12();
        Vector#(16, Struct26) x_29 = (update (x_27, (Bit#(4))'(4'hc),
        x_28));
        let x_30 <- rdResp_infoRam__00__13();
        Vector#(16, Struct26) x_31 = (update (x_29, (Bit#(4))'(4'hd),
        x_30));
        let x_32 <- rdResp_infoRam__00__14();
        Vector#(16, Struct26) x_33 = (update (x_31, (Bit#(4))'(4'he),
        x_32));
        let x_34 <- rdResp_infoRam__00__15();
        Vector#(16, Struct26) x_35 = (update (x_33, (Bit#(4))'(4'hf),
        x_34));
        Struct27 x_36 = (((((x_35)[(Bit#(4))'(4'h0)]).tag) == (x_1) ?
        (Struct27 {tm_hit : (Bool)'(True), tm_way : (Bit#(4))'(4'h0),
        tm_value : ((x_35)[(Bit#(4))'(4'h0)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h1)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h1), tm_value :
        ((x_35)[(Bit#(4))'(4'h1)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h2)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h2), tm_value :
        ((x_35)[(Bit#(4))'(4'h2)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h3)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h3), tm_value :
        ((x_35)[(Bit#(4))'(4'h3)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h4)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h4), tm_value :
        ((x_35)[(Bit#(4))'(4'h4)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h5)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h5), tm_value :
        ((x_35)[(Bit#(4))'(4'h5)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h6)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h6), tm_value :
        ((x_35)[(Bit#(4))'(4'h6)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h7)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h7), tm_value :
        ((x_35)[(Bit#(4))'(4'h7)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h8)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h8), tm_value :
        ((x_35)[(Bit#(4))'(4'h8)]).value}) :
        (((((x_35)[(Bit#(4))'(4'h9)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h9), tm_value :
        ((x_35)[(Bit#(4))'(4'h9)]).value}) :
        (((((x_35)[(Bit#(4))'(4'ha)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'ha), tm_value :
        ((x_35)[(Bit#(4))'(4'ha)]).value}) :
        (((((x_35)[(Bit#(4))'(4'hb)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hb), tm_value :
        ((x_35)[(Bit#(4))'(4'hb)]).value}) :
        (((((x_35)[(Bit#(4))'(4'hc)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hc), tm_value :
        ((x_35)[(Bit#(4))'(4'hc)]).value}) :
        (((((x_35)[(Bit#(4))'(4'hd)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hd), tm_value :
        ((x_35)[(Bit#(4))'(4'hd)]).value}) :
        (((((x_35)[(Bit#(4))'(4'he)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'he), tm_value :
        ((x_35)[(Bit#(4))'(4'he)]).value}) :
        (((((x_35)[(Bit#(4))'(4'hf)]).tag) == (x_1) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hf), tm_value :
        ((x_35)[(Bit#(4))'(4'hf)]).value}) :
        (unpack(0))))))))))))))))))))))))))))))))));
        Vector#(8, Struct28) x_37 = (unpack(0));
        let x_38 <- rdResp_edirRam__00__0();
        Vector#(8, Struct28) x_39 = (update (x_37, (Bit#(3))'(3'h0),
        x_38));
        let x_40 <- rdResp_edirRam__00__1();
        Vector#(8, Struct28) x_41 = (update (x_39, (Bit#(3))'(3'h1),
        x_40));
        let x_42 <- rdResp_edirRam__00__2();
        Vector#(8, Struct28) x_43 = (update (x_41, (Bit#(3))'(3'h2),
        x_42));
        let x_44 <- rdResp_edirRam__00__3();
        Vector#(8, Struct28) x_45 = (update (x_43, (Bit#(3))'(3'h3),
        x_44));
        let x_46 <- rdResp_edirRam__00__4();
        Vector#(8, Struct28) x_47 = (update (x_45, (Bit#(3))'(3'h4),
        x_46));
        let x_48 <- rdResp_edirRam__00__5();
        Vector#(8, Struct28) x_49 = (update (x_47, (Bit#(3))'(3'h5),
        x_48));
        let x_50 <- rdResp_edirRam__00__6();
        Vector#(8, Struct28) x_51 = (update (x_49, (Bit#(3))'(3'h6),
        x_50));
        let x_52 <- rdResp_edirRam__00__7();
        Vector#(8, Struct28) x_53 = (update (x_51, (Bit#(3))'(3'h7),
        x_52));
        Struct30 x_54 = (((((x_53)[(Bit#(3))'(3'h0)]).tag) == (x_1) ?
        (Struct30 {tm_hit : (Bool)'(True), tm_way : (Bit#(3))'(3'h0),
        tm_value : ((x_53)[(Bit#(3))'(3'h0)]).value}) :
        (((((x_53)[(Bit#(3))'(3'h1)]).tag) == (x_1) ? (Struct30 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h1), tm_value :
        ((x_53)[(Bit#(3))'(3'h1)]).value}) :
        (((((x_53)[(Bit#(3))'(3'h2)]).tag) == (x_1) ? (Struct30 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h2), tm_value :
        ((x_53)[(Bit#(3))'(3'h2)]).value}) :
        (((((x_53)[(Bit#(3))'(3'h3)]).tag) == (x_1) ? (Struct30 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h3), tm_value :
        ((x_53)[(Bit#(3))'(3'h3)]).value}) :
        (((((x_53)[(Bit#(3))'(3'h4)]).tag) == (x_1) ? (Struct30 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h4), tm_value :
        ((x_53)[(Bit#(3))'(3'h4)]).value}) :
        (((((x_53)[(Bit#(3))'(3'h5)]).tag) == (x_1) ? (Struct30 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h5), tm_value :
        ((x_53)[(Bit#(3))'(3'h5)]).value}) :
        (((((x_53)[(Bit#(3))'(3'h6)]).tag) == (x_1) ? (Struct30 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h6), tm_value :
        ((x_53)[(Bit#(3))'(3'h6)]).value}) :
        (((((x_53)[(Bit#(3))'(3'h7)]).tag) == (x_1) ? (Struct30 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h7), tm_value :
        ((x_53)[(Bit#(3))'(3'h7)]).value}) :
        (unpack(0))))))))))))))))));
        Struct29 x_55 = ((x_54).tm_value);
        Struct5 x_56 = ((! (((Bit#(3))'(3'h1)) <
        ((((x_53)[(Bit#(3))'(3'h0)]).value).mesi_edir_st)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((! (((Bit#(3))'(3'h1))
        < ((((x_53)[(Bit#(3))'(3'h1)]).value).mesi_edir_st)) ? (Struct5
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((!
        (((Bit#(3))'(3'h1)) <
        ((((x_53)[(Bit#(3))'(3'h2)]).value).mesi_edir_st)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((! (((Bit#(3))'(3'h1))
        < ((((x_53)[(Bit#(3))'(3'h3)]).value).mesi_edir_st)) ? (Struct5
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((!
        (((Bit#(3))'(3'h1)) <
        ((((x_53)[(Bit#(3))'(3'h4)]).value).mesi_edir_st)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((! (((Bit#(3))'(3'h1))
        < ((((x_53)[(Bit#(3))'(3'h5)]).value).mesi_edir_st)) ? (Struct5
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : ((!
        (((Bit#(3))'(3'h1)) <
        ((((x_53)[(Bit#(3))'(3'h6)]).value).mesi_edir_st)) ? (Struct5 {valid
        : (Bool)'(True), data : (Bit#(3))'(3'h6)}) : ((! (((Bit#(3))'(3'h1))
        < ((((x_53)[(Bit#(3))'(3'h7)]).value).mesi_edir_st)) ? (Struct5
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h7)}) : (Struct5 {valid :
        (Bool)'(False), data : unpack(0)})))))))))))))))));
        let x_57 <- repGetRs__00();
        Bit#(4) x_58 = (unpack(0));
        Bit#(8) x_59 = (unpack(0));
        Bit#(4) x_60 = ((! (((x_57)[(Bit#(4))'(4'hf)]) < (x_59)) ?
        ((Bit#(4))'(4'hf)) : (x_58)));
        Bit#(8) x_61 = ((! (((x_57)[(Bit#(4))'(4'hf)]) < (x_59)) ?
        ((x_57)[(Bit#(4))'(4'hf)]) : (x_59)));
        Bit#(4) x_62 = ((! (((x_57)[(Bit#(4))'(4'he)]) < (x_61)) ?
        ((Bit#(4))'(4'he)) : (x_60)));
        Bit#(8) x_63 = ((! (((x_57)[(Bit#(4))'(4'he)]) < (x_61)) ?
        ((x_57)[(Bit#(4))'(4'he)]) : (x_61)));
        Bit#(4) x_64 = ((! (((x_57)[(Bit#(4))'(4'hd)]) < (x_63)) ?
        ((Bit#(4))'(4'hd)) : (x_62)));
        Bit#(8) x_65 = ((! (((x_57)[(Bit#(4))'(4'hd)]) < (x_63)) ?
        ((x_57)[(Bit#(4))'(4'hd)]) : (x_63)));
        Bit#(4) x_66 = ((! (((x_57)[(Bit#(4))'(4'hc)]) < (x_65)) ?
        ((Bit#(4))'(4'hc)) : (x_64)));
        Bit#(8) x_67 = ((! (((x_57)[(Bit#(4))'(4'hc)]) < (x_65)) ?
        ((x_57)[(Bit#(4))'(4'hc)]) : (x_65)));
        Bit#(4) x_68 = ((! (((x_57)[(Bit#(4))'(4'hb)]) < (x_67)) ?
        ((Bit#(4))'(4'hb)) : (x_66)));
        Bit#(8) x_69 = ((! (((x_57)[(Bit#(4))'(4'hb)]) < (x_67)) ?
        ((x_57)[(Bit#(4))'(4'hb)]) : (x_67)));
        Bit#(4) x_70 = ((! (((x_57)[(Bit#(4))'(4'ha)]) < (x_69)) ?
        ((Bit#(4))'(4'ha)) : (x_68)));
        Bit#(8) x_71 = ((! (((x_57)[(Bit#(4))'(4'ha)]) < (x_69)) ?
        ((x_57)[(Bit#(4))'(4'ha)]) : (x_69)));
        Bit#(4) x_72 = ((! (((x_57)[(Bit#(4))'(4'h9)]) < (x_71)) ?
        ((Bit#(4))'(4'h9)) : (x_70)));
        Bit#(8) x_73 = ((! (((x_57)[(Bit#(4))'(4'h9)]) < (x_71)) ?
        ((x_57)[(Bit#(4))'(4'h9)]) : (x_71)));
        Bit#(4) x_74 = ((! (((x_57)[(Bit#(4))'(4'h8)]) < (x_73)) ?
        ((Bit#(4))'(4'h8)) : (x_72)));
        Bit#(8) x_75 = ((! (((x_57)[(Bit#(4))'(4'h8)]) < (x_73)) ?
        ((x_57)[(Bit#(4))'(4'h8)]) : (x_73)));
        Bit#(4) x_76 = ((! (((x_57)[(Bit#(4))'(4'h7)]) < (x_75)) ?
        ((Bit#(4))'(4'h7)) : (x_74)));
        Bit#(8) x_77 = ((! (((x_57)[(Bit#(4))'(4'h7)]) < (x_75)) ?
        ((x_57)[(Bit#(4))'(4'h7)]) : (x_75)));
        Bit#(4) x_78 = ((! (((x_57)[(Bit#(4))'(4'h6)]) < (x_77)) ?
        ((Bit#(4))'(4'h6)) : (x_76)));
        Bit#(8) x_79 = ((! (((x_57)[(Bit#(4))'(4'h6)]) < (x_77)) ?
        ((x_57)[(Bit#(4))'(4'h6)]) : (x_77)));
        Bit#(4) x_80 = ((! (((x_57)[(Bit#(4))'(4'h5)]) < (x_79)) ?
        ((Bit#(4))'(4'h5)) : (x_78)));
        Bit#(8) x_81 = ((! (((x_57)[(Bit#(4))'(4'h5)]) < (x_79)) ?
        ((x_57)[(Bit#(4))'(4'h5)]) : (x_79)));
        Bit#(4) x_82 = ((! (((x_57)[(Bit#(4))'(4'h4)]) < (x_81)) ?
        ((Bit#(4))'(4'h4)) : (x_80)));
        Bit#(8) x_83 = ((! (((x_57)[(Bit#(4))'(4'h4)]) < (x_81)) ?
        ((x_57)[(Bit#(4))'(4'h4)]) : (x_81)));
        Bit#(4) x_84 = ((! (((x_57)[(Bit#(4))'(4'h3)]) < (x_83)) ?
        ((Bit#(4))'(4'h3)) : (x_82)));
        Bit#(8) x_85 = ((! (((x_57)[(Bit#(4))'(4'h3)]) < (x_83)) ?
        ((x_57)[(Bit#(4))'(4'h3)]) : (x_83)));
        Bit#(4) x_86 = ((! (((x_57)[(Bit#(4))'(4'h2)]) < (x_85)) ?
        ((Bit#(4))'(4'h2)) : (x_84)));
        Bit#(8) x_87 = ((! (((x_57)[(Bit#(4))'(4'h2)]) < (x_85)) ?
        ((x_57)[(Bit#(4))'(4'h2)]) : (x_85)));
        Bit#(4) x_88 = ((! (((x_57)[(Bit#(4))'(4'h1)]) < (x_87)) ?
        ((Bit#(4))'(4'h1)) : (x_86)));
        Bit#(8) x_89 = ((! (((x_57)[(Bit#(4))'(4'h1)]) < (x_87)) ?
        ((x_57)[(Bit#(4))'(4'h1)]) : (x_87)));
        Bit#(4) x_90 = ((! (((x_57)[(Bit#(4))'(4'h0)]) < (x_89)) ?
        ((Bit#(4))'(4'h0)) : (x_88)));
        Bit#(8) x_91 = ((! (((x_57)[(Bit#(4))'(4'h0)]) < (x_89)) ?
        ((x_57)[(Bit#(4))'(4'h0)]) : (x_89)));
        when (! ((x_91) == ((Bit#(8))'(8'h0))), noAction);
        Struct26 x_92 = ((x_35)[x_90]);
        Bit#(50) x_93 = ((x_92).tag);
        Struct10 x_94 = ((x_92).value);
        Bit#(4) x_95 = (((x_36).tm_hit ? ((x_36).tm_way) : (x_90)));
        Struct9 x_96 = (Struct9 {info_index : x_2, info_hit : (x_36).tm_hit,
        info_way : x_95, edir_hit : (x_54).tm_hit, edir_way : (x_54).tm_way,
        edir_slot : x_56, info : ((x_36).tm_hit ? ((x_36).tm_value) :
        (Struct10 {mesi_owned : (x_55).mesi_edir_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : (x_55).mesi_edir_st, mesi_dir_sharers
        : (x_55).mesi_edir_sharers})), may_victim : Struct11 {mv_addr :
        {(x_93),({(x_2),((Bit#(5))'(5'h0))})}, mv_info : x_94}, reps :
        x_57});
        let x_97 <- rdReq_dataRam__00({(x_95),(x_2)});
        return x_96;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__00__valueRsLineRq
    (Struct17 x_0);
        let x_1 <- rdResp_dataRam__00();
        Bit#(64) x_2 = ((x_0).addr);
        Bit#(9) x_3 = ((x_2)[13:5]);
        Bit#(4) x_4 = ((x_0).info_way);
        Struct10 x_5 = ((x_0).info);
        Bool x_6 = ((! (((Bit#(3))'(3'h1)) < ((x_5).mesi_status))) && (!
        (((x_5).mesi_dir_st) == ((Bit#(3))'(3'h3)))));
        Struct5 x_7 = ((x_0).edir_slot);
        Bool x_8 = ((x_7).valid);
        Bit#(3) x_9 =
        ((x_7).data);
        if ((x_0).info_write)
            begin
            if ((((x_0).info_hit) || (! (x_6))) || (((! ((x_0).edir_hit)) &&
                (x_6)) && (! (x_8)))) begin
                Struct31 x_10 = (Struct31 {addr : x_3, datain : Struct26 {tag
                : (x_2)[63:14], value :
                x_5}});
                if ((x_4) == ((Bit#(4))'(4'h0))) begin
                    let x_11 <- wrReq_infoRam__00__0(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h1))) begin
                    let x_13 <- wrReq_infoRam__00__1(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h2))) begin
                    let x_15 <- wrReq_infoRam__00__2(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h3))) begin
                    let x_17 <- wrReq_infoRam__00__3(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h4))) begin
                    let x_19 <- wrReq_infoRam__00__4(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h5))) begin
                    let x_21 <- wrReq_infoRam__00__5(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h6))) begin
                    let x_23 <- wrReq_infoRam__00__6(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h7))) begin
                    let x_25 <- wrReq_infoRam__00__7(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h8))) begin
                    let x_27 <- wrReq_infoRam__00__8(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'h9))) begin
                    let x_29 <- wrReq_infoRam__00__9(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'ha))) begin
                    let x_31 <- wrReq_infoRam__00__10(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'hb))) begin
                    let x_33 <- wrReq_infoRam__00__11(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'hc))) begin
                    let x_35 <- wrReq_infoRam__00__12(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'hd))) begin
                    let x_37 <- wrReq_infoRam__00__13(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'he))) begin
                    let x_39 <- wrReq_infoRam__00__14(x_10);
                end else begin

                end
                if ((x_4) == ((Bit#(4))'(4'hf))) begin
                    let x_41 <- wrReq_infoRam__00__15(x_10);
                end else begin

                end
                if (! ((x_0).info_hit)) begin
                    Struct11 x_43 = ((x_0).may_victim);
                    Struct13 x_44 = (Struct13 {victim_valid : (Bool)'(True),
                    victim_addr : (x_43).mv_addr, victim_info :
                    (x_43).mv_info, victim_value : x_1, victim_req : Struct14
                    {valid : (Bool)'(False), data : unpack(0)}});
                    let x_45 <- victims__00__registerVictim(x_44);
                end else begin

                end
                let x_47 <- repAccess__00(Struct32 {acc_type : (!
                (((Bit#(3))'(3'h1)) < ((x_5).mesi_dir_st)) ?
                ((Bit#(1))'(1'h0)) : ((Bit#(1))'(1'h1))), acc_reps :
                (x_0).reps, acc_index : x_3, acc_way : x_4});
            end else begin

            end
            if (((! ((x_0).info_hit)) && (x_6)) && (((x_0).edir_hit) ||
                (x_8))) begin
                Bit#(3) x_49 = (((x_0).edir_hit ? ((x_0).edir_way) :
                (x_9)));
                Struct33 x_50 = (Struct33 {addr : (x_2)[13:5], datain :
                Struct28 {tag : (x_2)[63:14], value : Struct29
                {mesi_edir_owned : (x_5).mesi_owned, mesi_edir_st :
                (x_5).mesi_dir_st, mesi_edir_sharers :
                (x_5).mesi_dir_sharers}}});
                if ((x_49) == ((Bit#(3))'(3'h0))) begin
                    let x_51 <- wrReq_edirRam__00__0(x_50);
                end else begin

                end
                if ((x_49) == ((Bit#(3))'(3'h1))) begin
                    let x_53 <- wrReq_edirRam__00__1(x_50);
                end else begin

                end
                if ((x_49) == ((Bit#(3))'(3'h2))) begin
                    let x_55 <- wrReq_edirRam__00__2(x_50);
                end else begin

                end
                if ((x_49) == ((Bit#(3))'(3'h3))) begin
                    let x_57 <- wrReq_edirRam__00__3(x_50);
                end else begin

                end
                if ((x_49) == ((Bit#(3))'(3'h4))) begin
                    let x_59 <- wrReq_edirRam__00__4(x_50);
                end else begin

                end
                if ((x_49) == ((Bit#(3))'(3'h5))) begin
                    let x_61 <- wrReq_edirRam__00__5(x_50);
                end else begin

                end
                if ((x_49) == ((Bit#(3))'(3'h6))) begin
                    let x_63 <- wrReq_edirRam__00__6(x_50);
                end else begin

                end
                if ((x_49) == ((Bit#(3))'(3'h7))) begin
                    let x_65 <- wrReq_edirRam__00__7(x_50);
                end else begin

                end
            end else
                begin
                if ((x_0).edir_hit) begin
                    Bit#(3) x_67 = ((x_0).edir_way);
                    Struct33 x_68 = (Struct33 {addr : (x_2)[13:5], datain :
                    Struct28 {tag : (x_2)[63:14], value : Struct29
                    {mesi_edir_owned : (x_5).mesi_owned, mesi_edir_st :
                    (x_5).mesi_dir_st, mesi_edir_sharers :
                    (x_5).mesi_dir_sharers}}});
                    if ((x_67) == ((Bit#(3))'(3'h0))) begin
                        let x_69 <- wrReq_edirRam__00__0(x_68);
                    end else begin

                    end
                    if ((x_67) == ((Bit#(3))'(3'h1))) begin
                        let x_71 <- wrReq_edirRam__00__1(x_68);
                    end else begin

                    end
                    if ((x_67) == ((Bit#(3))'(3'h2))) begin
                        let x_73 <- wrReq_edirRam__00__2(x_68);
                    end else begin

                    end
                    if ((x_67) == ((Bit#(3))'(3'h3))) begin
                        let x_75 <- wrReq_edirRam__00__3(x_68);
                    end else begin

                    end
                    if ((x_67) == ((Bit#(3))'(3'h4))) begin
                        let x_77 <- wrReq_edirRam__00__4(x_68);
                    end else begin

                    end
                    if ((x_67) == ((Bit#(3))'(3'h5))) begin
                        let x_79 <- wrReq_edirRam__00__5(x_68);
                    end else begin

                    end
                    if ((x_67) == ((Bit#(3))'(3'h6))) begin
                        let x_81 <- wrReq_edirRam__00__6(x_68);
                    end else begin

                    end
                    if ((x_67) == ((Bit#(3))'(3'h7))) begin
                        let x_83 <- wrReq_edirRam__00__7(x_68);
                    end else begin

                    end
                end else begin

                end
            end
        end else begin

        end
        if ((x_0).value_write) begin
            Struct34 x_88 = (Struct34 {addr : {(x_4),((x_2)[13:5])}, datain :
            (x_0).value});
            let x_89 <- wrReq_dataRam__00(x_88);
        end else begin

        end
        return x_1;
    endmethod
endmodule

interface Module129;
    method Action cache__000__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct41) cache__000__infoRsValueRq (Bit#(64) x_0);
    method ActionValue#(Vector#(4, Bit#(64))) cache__000__valueRsLineRq
    (Struct46 x_0);
endinterface

module mkModule129#(function Action wrReq_dataRam__000(Struct54 _),
    function Action repAccess__000(Struct53 _),
    function Action victims__000__registerVictim(Struct44 _),
    function Action wrReq_infoRam__000__3(Struct52 _),
    function Action wrReq_infoRam__000__2(Struct52 _),
    function Action wrReq_infoRam__000__1(Struct52 _),
    function Action wrReq_infoRam__000__0(Struct52 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__000(),
    function Action rdReq_dataRam__000(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__000(),
    function ActionValue#(Struct50) rdResp_infoRam__000__3(),
    function ActionValue#(Struct50) rdResp_infoRam__000__2(),
    function ActionValue#(Struct50) rdResp_infoRam__000__1(),
    function ActionValue#(Struct50) rdResp_infoRam__000__0(),
    function Action repGetRq__000(Bit#(8) _),
    function Action rdReq_infoRam__000__3(Bit#(8) _),
    function Action rdReq_infoRam__000__2(Bit#(8) _),
    function Action rdReq_infoRam__000__1(Bit#(8) _),
    function Action rdReq_infoRam__000__0(Bit#(8) _))
    (Module129);

    // No rules in this module

    method Action cache__000__infoRq (Bit#(64) x_0);
        Bit#(8) x_1 = ((x_0)[12:5]);
        let x_2 <- rdReq_infoRam__000__0(x_1);
        let x_3 <- rdReq_infoRam__000__1(x_1);
        let x_4 <- rdReq_infoRam__000__2(x_1);
        let x_5 <- rdReq_infoRam__000__3(x_1);
        let x_6 <- repGetRq__000(x_1);
    endmethod

    method ActionValue#(Struct41) cache__000__infoRsValueRq (Bit#(64) x_0);
        Bit#(51) x_1 = ((x_0)[63:13]);
        Bit#(8) x_2 = ((x_0)[12:5]);
        Vector#(4, Struct50) x_3 = (unpack(0));
        let x_4 <- rdResp_infoRam__000__0();
        Vector#(4, Struct50) x_5 = (update (x_3, (Bit#(2))'(2'h0), x_4));
        let x_6 <- rdResp_infoRam__000__1();
        Vector#(4, Struct50) x_7 = (update (x_5, (Bit#(2))'(2'h1), x_6));
        let x_8 <- rdResp_infoRam__000__2();
        Vector#(4, Struct50) x_9 = (update (x_7, (Bit#(2))'(2'h2), x_8));
        let x_10 <- rdResp_infoRam__000__3();
        Vector#(4, Struct50) x_11 = (update (x_9, (Bit#(2))'(2'h3),
        x_10));
        Struct51 x_12 = (((((x_11)[(Bit#(2))'(2'h0)]).tag) == (x_1) ?
        (Struct51 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_11)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h1)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_11)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h2)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_11)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h3)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_11)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
        let x_13 <- repGetRs__000();
        Bit#(2) x_14 = (unpack(0));
        Bit#(8) x_15 = (unpack(0));
        Bit#(2) x_16 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((Bit#(2))'(2'h3)) : (x_14)));
        Bit#(8) x_17 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((x_13)[(Bit#(2))'(2'h3)]) : (x_15)));
        Bit#(2) x_18 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((Bit#(2))'(2'h2)) : (x_16)));
        Bit#(8) x_19 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((x_13)[(Bit#(2))'(2'h2)]) : (x_17)));
        Bit#(2) x_20 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((Bit#(2))'(2'h1)) : (x_18)));
        Bit#(8) x_21 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((x_13)[(Bit#(2))'(2'h1)]) : (x_19)));
        Bit#(2) x_22 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((Bit#(2))'(2'h0)) : (x_20)));
        Bit#(8) x_23 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((x_13)[(Bit#(2))'(2'h0)]) : (x_21)));
        when (! ((x_23) == ((Bit#(8))'(8'h0))), noAction);
        Struct50 x_24 = ((x_11)[x_22]);
        Bit#(51) x_25 = ((x_24).tag);
        Struct10 x_26 = ((x_24).value);
        Bit#(2) x_27 = (((x_12).tm_hit ? ((x_12).tm_way) : (x_22)));
        Struct41 x_28 = (Struct41 {info_index : x_2, info_hit :
        (x_12).tm_hit, info_way : x_27, edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_12).tm_value, may_victim
        : Struct11 {mv_addr : {(x_25),({(x_2),((Bit#(5))'(5'h0))})}, mv_info
        : x_26}, reps : x_13});
        let x_29 <- rdReq_dataRam__000({(x_27),(x_2)});
        return x_28;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__000__valueRsLineRq
    (Struct46 x_0);
        let x_1 <- rdResp_dataRam__000();
        Bit#(64) x_2 = ((x_0).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Bit#(2) x_4 = ((x_0).info_way);
        Struct10 x_5 =
        ((x_0).info);
        if ((x_0).info_write) begin
            Struct52 x_6 = (Struct52 {addr : x_3, datain : Struct50 {tag :
            (x_2)[63:13], value :
            x_5}});
            if ((x_4) == ((Bit#(2))'(2'h0))) begin
                let x_7 <- wrReq_infoRam__000__0(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h1))) begin
                let x_9 <- wrReq_infoRam__000__1(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h2))) begin
                let x_11 <- wrReq_infoRam__000__2(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h3))) begin
                let x_13 <- wrReq_infoRam__000__3(x_6);
            end else begin

            end
            if (! ((x_0).info_hit)) begin
                Struct11 x_15 = ((x_0).may_victim);
                Struct44 x_16 = (Struct44 {victim_valid : (Bool)'(True),
                victim_addr : (x_15).mv_addr, victim_info : (x_15).mv_info,
                victim_value : x_1, victim_req : Struct5 {valid :
                (Bool)'(False), data : unpack(0)}});
                let x_17 <- victims__000__registerVictim(x_16);
            end else begin

            end
            let x_19 <- repAccess__000(Struct53 {acc_type : (!
            (((Bit#(3))'(3'h1)) < ((x_5).mesi_dir_st)) ? ((Bit#(1))'(1'h0)) :
            ((Bit#(1))'(1'h1))), acc_reps : (x_0).reps, acc_index : x_3,
            acc_way : x_4});
        end else begin

        end
        if ((x_0).value_write) begin
            Struct54 x_21 = (Struct54 {addr : {(x_4),((x_2)[12:5])}, datain :
            (x_0).value});
            let x_22 <- wrReq_dataRam__000(x_21);
        end else begin

        end
        return x_1;
    endmethod
endmodule

interface Module130;
    method Action cache__001__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct41) cache__001__infoRsValueRq (Bit#(64) x_0);
    method ActionValue#(Vector#(4, Bit#(64))) cache__001__valueRsLineRq
    (Struct46 x_0);
endinterface

module mkModule130#(function Action wrReq_dataRam__001(Struct54 _),
    function Action repAccess__001(Struct53 _),
    function Action victims__001__registerVictim(Struct44 _),
    function Action wrReq_infoRam__001__3(Struct52 _),
    function Action wrReq_infoRam__001__2(Struct52 _),
    function Action wrReq_infoRam__001__1(Struct52 _),
    function Action wrReq_infoRam__001__0(Struct52 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__001(),
    function Action rdReq_dataRam__001(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__001(),
    function ActionValue#(Struct50) rdResp_infoRam__001__3(),
    function ActionValue#(Struct50) rdResp_infoRam__001__2(),
    function ActionValue#(Struct50) rdResp_infoRam__001__1(),
    function ActionValue#(Struct50) rdResp_infoRam__001__0(),
    function Action repGetRq__001(Bit#(8) _),
    function Action rdReq_infoRam__001__3(Bit#(8) _),
    function Action rdReq_infoRam__001__2(Bit#(8) _),
    function Action rdReq_infoRam__001__1(Bit#(8) _),
    function Action rdReq_infoRam__001__0(Bit#(8) _))
    (Module130);

    // No rules in this module

    method Action cache__001__infoRq (Bit#(64) x_0);
        Bit#(8) x_1 = ((x_0)[12:5]);
        let x_2 <- rdReq_infoRam__001__0(x_1);
        let x_3 <- rdReq_infoRam__001__1(x_1);
        let x_4 <- rdReq_infoRam__001__2(x_1);
        let x_5 <- rdReq_infoRam__001__3(x_1);
        let x_6 <- repGetRq__001(x_1);
    endmethod

    method ActionValue#(Struct41) cache__001__infoRsValueRq (Bit#(64) x_0);
        Bit#(51) x_1 = ((x_0)[63:13]);
        Bit#(8) x_2 = ((x_0)[12:5]);
        Vector#(4, Struct50) x_3 = (unpack(0));
        let x_4 <- rdResp_infoRam__001__0();
        Vector#(4, Struct50) x_5 = (update (x_3, (Bit#(2))'(2'h0), x_4));
        let x_6 <- rdResp_infoRam__001__1();
        Vector#(4, Struct50) x_7 = (update (x_5, (Bit#(2))'(2'h1), x_6));
        let x_8 <- rdResp_infoRam__001__2();
        Vector#(4, Struct50) x_9 = (update (x_7, (Bit#(2))'(2'h2), x_8));
        let x_10 <- rdResp_infoRam__001__3();
        Vector#(4, Struct50) x_11 = (update (x_9, (Bit#(2))'(2'h3),
        x_10));
        Struct51 x_12 = (((((x_11)[(Bit#(2))'(2'h0)]).tag) == (x_1) ?
        (Struct51 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_11)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h1)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_11)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h2)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_11)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h3)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_11)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
        let x_13 <- repGetRs__001();
        Bit#(2) x_14 = (unpack(0));
        Bit#(8) x_15 = (unpack(0));
        Bit#(2) x_16 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((Bit#(2))'(2'h3)) : (x_14)));
        Bit#(8) x_17 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((x_13)[(Bit#(2))'(2'h3)]) : (x_15)));
        Bit#(2) x_18 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((Bit#(2))'(2'h2)) : (x_16)));
        Bit#(8) x_19 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((x_13)[(Bit#(2))'(2'h2)]) : (x_17)));
        Bit#(2) x_20 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((Bit#(2))'(2'h1)) : (x_18)));
        Bit#(8) x_21 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((x_13)[(Bit#(2))'(2'h1)]) : (x_19)));
        Bit#(2) x_22 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((Bit#(2))'(2'h0)) : (x_20)));
        Bit#(8) x_23 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((x_13)[(Bit#(2))'(2'h0)]) : (x_21)));
        when (! ((x_23) == ((Bit#(8))'(8'h0))), noAction);
        Struct50 x_24 = ((x_11)[x_22]);
        Bit#(51) x_25 = ((x_24).tag);
        Struct10 x_26 = ((x_24).value);
        Bit#(2) x_27 = (((x_12).tm_hit ? ((x_12).tm_way) : (x_22)));
        Struct41 x_28 = (Struct41 {info_index : x_2, info_hit :
        (x_12).tm_hit, info_way : x_27, edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_12).tm_value, may_victim
        : Struct11 {mv_addr : {(x_25),({(x_2),((Bit#(5))'(5'h0))})}, mv_info
        : x_26}, reps : x_13});
        let x_29 <- rdReq_dataRam__001({(x_27),(x_2)});
        return x_28;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__001__valueRsLineRq
    (Struct46 x_0);
        let x_1 <- rdResp_dataRam__001();
        Bit#(64) x_2 = ((x_0).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Bit#(2) x_4 = ((x_0).info_way);
        Struct10 x_5 =
        ((x_0).info);
        if ((x_0).info_write) begin
            Struct52 x_6 = (Struct52 {addr : x_3, datain : Struct50 {tag :
            (x_2)[63:13], value :
            x_5}});
            if ((x_4) == ((Bit#(2))'(2'h0))) begin
                let x_7 <- wrReq_infoRam__001__0(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h1))) begin
                let x_9 <- wrReq_infoRam__001__1(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h2))) begin
                let x_11 <- wrReq_infoRam__001__2(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h3))) begin
                let x_13 <- wrReq_infoRam__001__3(x_6);
            end else begin

            end
            if (! ((x_0).info_hit)) begin
                Struct11 x_15 = ((x_0).may_victim);
                Struct44 x_16 = (Struct44 {victim_valid : (Bool)'(True),
                victim_addr : (x_15).mv_addr, victim_info : (x_15).mv_info,
                victim_value : x_1, victim_req : Struct5 {valid :
                (Bool)'(False), data : unpack(0)}});
                let x_17 <- victims__001__registerVictim(x_16);
            end else begin

            end
            let x_19 <- repAccess__001(Struct53 {acc_type : (!
            (((Bit#(3))'(3'h1)) < ((x_5).mesi_dir_st)) ? ((Bit#(1))'(1'h0)) :
            ((Bit#(1))'(1'h1))), acc_reps : (x_0).reps, acc_index : x_3,
            acc_way : x_4});
        end else begin

        end
        if ((x_0).value_write) begin
            Struct54 x_21 = (Struct54 {addr : {(x_4),((x_2)[12:5])}, datain :
            (x_0).value});
            let x_22 <- wrReq_dataRam__001(x_21);
        end else begin

        end
        return x_1;
    endmethod
endmodule

interface Module131;
    method Action cache__002__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct41) cache__002__infoRsValueRq (Bit#(64) x_0);
    method ActionValue#(Vector#(4, Bit#(64))) cache__002__valueRsLineRq
    (Struct46 x_0);
endinterface

module mkModule131#(function Action wrReq_dataRam__002(Struct54 _),
    function Action repAccess__002(Struct53 _),
    function Action victims__002__registerVictim(Struct44 _),
    function Action wrReq_infoRam__002__3(Struct52 _),
    function Action wrReq_infoRam__002__2(Struct52 _),
    function Action wrReq_infoRam__002__1(Struct52 _),
    function Action wrReq_infoRam__002__0(Struct52 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__002(),
    function Action rdReq_dataRam__002(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__002(),
    function ActionValue#(Struct50) rdResp_infoRam__002__3(),
    function ActionValue#(Struct50) rdResp_infoRam__002__2(),
    function ActionValue#(Struct50) rdResp_infoRam__002__1(),
    function ActionValue#(Struct50) rdResp_infoRam__002__0(),
    function Action repGetRq__002(Bit#(8) _),
    function Action rdReq_infoRam__002__3(Bit#(8) _),
    function Action rdReq_infoRam__002__2(Bit#(8) _),
    function Action rdReq_infoRam__002__1(Bit#(8) _),
    function Action rdReq_infoRam__002__0(Bit#(8) _))
    (Module131);

    // No rules in this module

    method Action cache__002__infoRq (Bit#(64) x_0);
        Bit#(8) x_1 = ((x_0)[12:5]);
        let x_2 <- rdReq_infoRam__002__0(x_1);
        let x_3 <- rdReq_infoRam__002__1(x_1);
        let x_4 <- rdReq_infoRam__002__2(x_1);
        let x_5 <- rdReq_infoRam__002__3(x_1);
        let x_6 <- repGetRq__002(x_1);
    endmethod

    method ActionValue#(Struct41) cache__002__infoRsValueRq (Bit#(64) x_0);
        Bit#(51) x_1 = ((x_0)[63:13]);
        Bit#(8) x_2 = ((x_0)[12:5]);
        Vector#(4, Struct50) x_3 = (unpack(0));
        let x_4 <- rdResp_infoRam__002__0();
        Vector#(4, Struct50) x_5 = (update (x_3, (Bit#(2))'(2'h0), x_4));
        let x_6 <- rdResp_infoRam__002__1();
        Vector#(4, Struct50) x_7 = (update (x_5, (Bit#(2))'(2'h1), x_6));
        let x_8 <- rdResp_infoRam__002__2();
        Vector#(4, Struct50) x_9 = (update (x_7, (Bit#(2))'(2'h2), x_8));
        let x_10 <- rdResp_infoRam__002__3();
        Vector#(4, Struct50) x_11 = (update (x_9, (Bit#(2))'(2'h3),
        x_10));
        Struct51 x_12 = (((((x_11)[(Bit#(2))'(2'h0)]).tag) == (x_1) ?
        (Struct51 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_11)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h1)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_11)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h2)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_11)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h3)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_11)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
        let x_13 <- repGetRs__002();
        Bit#(2) x_14 = (unpack(0));
        Bit#(8) x_15 = (unpack(0));
        Bit#(2) x_16 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((Bit#(2))'(2'h3)) : (x_14)));
        Bit#(8) x_17 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((x_13)[(Bit#(2))'(2'h3)]) : (x_15)));
        Bit#(2) x_18 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((Bit#(2))'(2'h2)) : (x_16)));
        Bit#(8) x_19 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((x_13)[(Bit#(2))'(2'h2)]) : (x_17)));
        Bit#(2) x_20 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((Bit#(2))'(2'h1)) : (x_18)));
        Bit#(8) x_21 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((x_13)[(Bit#(2))'(2'h1)]) : (x_19)));
        Bit#(2) x_22 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((Bit#(2))'(2'h0)) : (x_20)));
        Bit#(8) x_23 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((x_13)[(Bit#(2))'(2'h0)]) : (x_21)));
        when (! ((x_23) == ((Bit#(8))'(8'h0))), noAction);
        Struct50 x_24 = ((x_11)[x_22]);
        Bit#(51) x_25 = ((x_24).tag);
        Struct10 x_26 = ((x_24).value);
        Bit#(2) x_27 = (((x_12).tm_hit ? ((x_12).tm_way) : (x_22)));
        Struct41 x_28 = (Struct41 {info_index : x_2, info_hit :
        (x_12).tm_hit, info_way : x_27, edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_12).tm_value, may_victim
        : Struct11 {mv_addr : {(x_25),({(x_2),((Bit#(5))'(5'h0))})}, mv_info
        : x_26}, reps : x_13});
        let x_29 <- rdReq_dataRam__002({(x_27),(x_2)});
        return x_28;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__002__valueRsLineRq
    (Struct46 x_0);
        let x_1 <- rdResp_dataRam__002();
        Bit#(64) x_2 = ((x_0).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Bit#(2) x_4 = ((x_0).info_way);
        Struct10 x_5 =
        ((x_0).info);
        if ((x_0).info_write) begin
            Struct52 x_6 = (Struct52 {addr : x_3, datain : Struct50 {tag :
            (x_2)[63:13], value :
            x_5}});
            if ((x_4) == ((Bit#(2))'(2'h0))) begin
                let x_7 <- wrReq_infoRam__002__0(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h1))) begin
                let x_9 <- wrReq_infoRam__002__1(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h2))) begin
                let x_11 <- wrReq_infoRam__002__2(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h3))) begin
                let x_13 <- wrReq_infoRam__002__3(x_6);
            end else begin

            end
            if (! ((x_0).info_hit)) begin
                Struct11 x_15 = ((x_0).may_victim);
                Struct44 x_16 = (Struct44 {victim_valid : (Bool)'(True),
                victim_addr : (x_15).mv_addr, victim_info : (x_15).mv_info,
                victim_value : x_1, victim_req : Struct5 {valid :
                (Bool)'(False), data : unpack(0)}});
                let x_17 <- victims__002__registerVictim(x_16);
            end else begin

            end
            let x_19 <- repAccess__002(Struct53 {acc_type : (!
            (((Bit#(3))'(3'h1)) < ((x_5).mesi_dir_st)) ? ((Bit#(1))'(1'h0)) :
            ((Bit#(1))'(1'h1))), acc_reps : (x_0).reps, acc_index : x_3,
            acc_way : x_4});
        end else begin

        end
        if ((x_0).value_write) begin
            Struct54 x_21 = (Struct54 {addr : {(x_4),((x_2)[12:5])}, datain :
            (x_0).value});
            let x_22 <- wrReq_dataRam__002(x_21);
        end else begin

        end
        return x_1;
    endmethod
endmodule

interface Module132;
    method Action cache__003__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct41) cache__003__infoRsValueRq (Bit#(64) x_0);
    method ActionValue#(Vector#(4, Bit#(64))) cache__003__valueRsLineRq
    (Struct46 x_0);
endinterface

module mkModule132#(function Action wrReq_dataRam__003(Struct54 _),
    function Action repAccess__003(Struct53 _),
    function Action victims__003__registerVictim(Struct44 _),
    function Action wrReq_infoRam__003__3(Struct52 _),
    function Action wrReq_infoRam__003__2(Struct52 _),
    function Action wrReq_infoRam__003__1(Struct52 _),
    function Action wrReq_infoRam__003__0(Struct52 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__003(),
    function Action rdReq_dataRam__003(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__003(),
    function ActionValue#(Struct50) rdResp_infoRam__003__3(),
    function ActionValue#(Struct50) rdResp_infoRam__003__2(),
    function ActionValue#(Struct50) rdResp_infoRam__003__1(),
    function ActionValue#(Struct50) rdResp_infoRam__003__0(),
    function Action repGetRq__003(Bit#(8) _),
    function Action rdReq_infoRam__003__3(Bit#(8) _),
    function Action rdReq_infoRam__003__2(Bit#(8) _),
    function Action rdReq_infoRam__003__1(Bit#(8) _),
    function Action rdReq_infoRam__003__0(Bit#(8) _))
    (Module132);

    // No rules in this module

    method Action cache__003__infoRq (Bit#(64) x_0);
        Bit#(8) x_1 = ((x_0)[12:5]);
        let x_2 <- rdReq_infoRam__003__0(x_1);
        let x_3 <- rdReq_infoRam__003__1(x_1);
        let x_4 <- rdReq_infoRam__003__2(x_1);
        let x_5 <- rdReq_infoRam__003__3(x_1);
        let x_6 <- repGetRq__003(x_1);
    endmethod

    method ActionValue#(Struct41) cache__003__infoRsValueRq (Bit#(64) x_0);
        Bit#(51) x_1 = ((x_0)[63:13]);
        Bit#(8) x_2 = ((x_0)[12:5]);
        Vector#(4, Struct50) x_3 = (unpack(0));
        let x_4 <- rdResp_infoRam__003__0();
        Vector#(4, Struct50) x_5 = (update (x_3, (Bit#(2))'(2'h0), x_4));
        let x_6 <- rdResp_infoRam__003__1();
        Vector#(4, Struct50) x_7 = (update (x_5, (Bit#(2))'(2'h1), x_6));
        let x_8 <- rdResp_infoRam__003__2();
        Vector#(4, Struct50) x_9 = (update (x_7, (Bit#(2))'(2'h2), x_8));
        let x_10 <- rdResp_infoRam__003__3();
        Vector#(4, Struct50) x_11 = (update (x_9, (Bit#(2))'(2'h3),
        x_10));
        Struct51 x_12 = (((((x_11)[(Bit#(2))'(2'h0)]).tag) == (x_1) ?
        (Struct51 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_11)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h1)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_11)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h2)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_11)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_11)[(Bit#(2))'(2'h3)]).tag) == (x_1) ? (Struct51 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_11)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
        let x_13 <- repGetRs__003();
        Bit#(2) x_14 = (unpack(0));
        Bit#(8) x_15 = (unpack(0));
        Bit#(2) x_16 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((Bit#(2))'(2'h3)) : (x_14)));
        Bit#(8) x_17 = ((! (((x_13)[(Bit#(2))'(2'h3)]) < (x_15)) ?
        ((x_13)[(Bit#(2))'(2'h3)]) : (x_15)));
        Bit#(2) x_18 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((Bit#(2))'(2'h2)) : (x_16)));
        Bit#(8) x_19 = ((! (((x_13)[(Bit#(2))'(2'h2)]) < (x_17)) ?
        ((x_13)[(Bit#(2))'(2'h2)]) : (x_17)));
        Bit#(2) x_20 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((Bit#(2))'(2'h1)) : (x_18)));
        Bit#(8) x_21 = ((! (((x_13)[(Bit#(2))'(2'h1)]) < (x_19)) ?
        ((x_13)[(Bit#(2))'(2'h1)]) : (x_19)));
        Bit#(2) x_22 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((Bit#(2))'(2'h0)) : (x_20)));
        Bit#(8) x_23 = ((! (((x_13)[(Bit#(2))'(2'h0)]) < (x_21)) ?
        ((x_13)[(Bit#(2))'(2'h0)]) : (x_21)));
        when (! ((x_23) == ((Bit#(8))'(8'h0))), noAction);
        Struct50 x_24 = ((x_11)[x_22]);
        Bit#(51) x_25 = ((x_24).tag);
        Struct10 x_26 = ((x_24).value);
        Bit#(2) x_27 = (((x_12).tm_hit ? ((x_12).tm_way) : (x_22)));
        Struct41 x_28 = (Struct41 {info_index : x_2, info_hit :
        (x_12).tm_hit, info_way : x_27, edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_12).tm_value, may_victim
        : Struct11 {mv_addr : {(x_25),({(x_2),((Bit#(5))'(5'h0))})}, mv_info
        : x_26}, reps : x_13});
        let x_29 <- rdReq_dataRam__003({(x_27),(x_2)});
        return x_28;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__003__valueRsLineRq
    (Struct46 x_0);
        let x_1 <- rdResp_dataRam__003();
        Bit#(64) x_2 = ((x_0).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Bit#(2) x_4 = ((x_0).info_way);
        Struct10 x_5 =
        ((x_0).info);
        if ((x_0).info_write) begin
            Struct52 x_6 = (Struct52 {addr : x_3, datain : Struct50 {tag :
            (x_2)[63:13], value :
            x_5}});
            if ((x_4) == ((Bit#(2))'(2'h0))) begin
                let x_7 <- wrReq_infoRam__003__0(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h1))) begin
                let x_9 <- wrReq_infoRam__003__1(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h2))) begin
                let x_11 <- wrReq_infoRam__003__2(x_6);
            end else begin

            end
            if ((x_4) == ((Bit#(2))'(2'h3))) begin
                let x_13 <- wrReq_infoRam__003__3(x_6);
            end else begin

            end
            if (! ((x_0).info_hit)) begin
                Struct11 x_15 = ((x_0).may_victim);
                Struct44 x_16 = (Struct44 {victim_valid : (Bool)'(True),
                victim_addr : (x_15).mv_addr, victim_info : (x_15).mv_info,
                victim_value : x_1, victim_req : Struct5 {valid :
                (Bool)'(False), data : unpack(0)}});
                let x_17 <- victims__003__registerVictim(x_16);
            end else begin

            end
            let x_19 <- repAccess__003(Struct53 {acc_type : (!
            (((Bit#(3))'(3'h1)) < ((x_5).mesi_dir_st)) ? ((Bit#(1))'(1'h0)) :
            ((Bit#(1))'(1'h1))), acc_reps : (x_0).reps, acc_index : x_3,
            acc_way : x_4});
        end else begin

        end
        if ((x_0).value_write) begin
            Struct54 x_21 = (Struct54 {addr : {(x_4),((x_2)[12:5])}, datain :
            (x_0).value});
            let x_22 <- wrReq_dataRam__003(x_21);
        end else begin

        end
        return x_1;
    endmethod
endmodule

interface Module133;

endinterface

module mkModule133#(function Action canImm_00(Bit#(64) _),
    function Action victims__00__setVictimRq(Struct25 _),
    function ActionValue#(Bit#(4)) setULImm_00(Struct1 _),
    function ActionValue#(Struct13) victims__00__getFirstVictim(),
    function Action transferUpDown_00(Struct24 _),
    function Action broadcast_parentChildren00(Struct22 _),
    function Action registerDL_00(Struct21 _),
    function Action registerUL_00(Struct20 _),
    function Action makeEnq_parentChildren00(Struct19 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__00__valueRsLineRq(Struct17 _),
    function Action victims__00__setVictim(Struct18 _),
    function ActionValue#(Struct15) getMSHR_00(Bit#(4) _),
    function ActionValue#(Struct12) deq_fifoL2E_00(),
    function ActionValue#(Struct13) victims__00__getVictim(Bit#(3) _),
    function Action enq_fifoL2E_00(Struct12 _),
    function ActionValue#(Struct9) cache__00__infoRsValueRq(Bit#(64) _),
    function ActionValue#(Struct6) deq_fifoI2L_00(),
    function Action enq_fifoI2L_00(Struct6 _),
    function Action cache__00__infoRq(Bit#(64) _),
    function ActionValue#(Struct6) deq_fifoN2I_00(),
    function ActionValue#(Struct8) getDLReady_00(),
    function Action addRs_00(Struct7 _),
    function ActionValue#(Struct2) deq_fifoCRsInput_00(),
    function ActionValue#(Struct4) getCRqSlot_00(Struct3 _),
    function ActionValue#(Bool) victims__00__hasVictim(),
    function ActionValue#(Struct2) deq_fifoCRqInput_00(),
    function Action releaseMSHR_00(Bit#(4) _),
    function ActionValue#(Bit#(4)) victims__00__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct3) getWait_00(),
    function Action startRelease_00(Bit#(4) _),
    function ActionValue#(Bit#(4)) getULReady_00(Bit#(64) _),
    function Action enq_fifoN2I_00(Struct6 _),
    function ActionValue#(Struct5) victims__00__findVictim(Bit#(64) _),
    function ActionValue#(Struct4) getPRqSlot_00(Struct3 _),
    function ActionValue#(Struct2) deq_fifoPInput_00())
    (Module133);

    rule rule_in_prq_00;
        $display ("Rule fired: rule_in_prq_00 at %t", $time);
        let x_0 <- deq_fifoPInput_00();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_00(Struct3 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).in_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- victims__00__findVictim((x_2).addr);
            Struct6 x_5 = (Struct6 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id,
            ir_by_victim : x_4});
            let x_6 <- enq_fifoN2I_00(x_5);
        end else begin

        end
    endrule

    rule rule_in_prs_00;
        $display ("Rule fired: rule_in_prs_00 at %t", $time);
        let x_0 <- deq_fifoPInput_00();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- getULReady_00((x_2).addr);
        let x_4 <- startRelease_00(x_3);
        let x_5 <- victims__00__findVictim((x_2).addr);
        Struct6 x_6 = (Struct6 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : x_3, ir_by_victim :
        x_5});
        let x_7 <- enq_fifoN2I_00(x_6);
    endrule

    rule rule_in_retry_00;
        $display ("Rule fired: rule_in_retry_00 at %t", $time);
        let x_0 <- getWait_00();
        Struct1 x_1 = ((x_0).r_msg);
        let x_2 <- victims__00__findVictim((x_1).addr);
        Struct6 x_3 = (Struct6 {ir_is_rs_rel : (Bool)'(False), ir_msg : x_1,
        ir_msg_from : (x_0).r_msg_from, ir_mshr_id : (x_0).r_id, ir_by_victim
        : x_2});
        let x_4 <- enq_fifoN2I_00(x_3);
    endrule

    rule rule_in_invrs_00;
        $display ("Rule fired: rule_in_invrs_00 at %t", $time);
        let x_0 <- deq_fifoPInput_00();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- getULReady_00((x_2).addr);
        let x_4 <- victims__00__releaseVictim((x_2).addr);
        let x_5 <- releaseMSHR_00(x_3);
    endrule

    rule rule_in_crq_00;
        $display ("Rule fired: rule_in_crq_00 at %t", $time);
        let x_0 <- deq_fifoCRqInput_00();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when (((x_1)[3:2]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- victims__00__hasVictim();
        when (! (x_3), noAction);
        let x_4 <- getCRqSlot_00(Struct3 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_4).s_has_slot,
        noAction);
        if (! ((x_4).s_conflict)) begin
            let x_5 <- victims__00__findVictim((x_2).addr);
            Struct6 x_6 = (Struct6 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_4).s_id,
            ir_by_victim : x_5});
            let x_7 <- enq_fifoN2I_00(x_6);
        end else begin

        end
    endrule

    rule rule_in_crs_00;
        $display ("Rule fired: rule_in_crs_00 at %t", $time);
        let x_0 <- deq_fifoCRsInput_00();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when (((x_1)[3:2]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_00(Struct7 {r_midx : (x_1)[1:0], r_msg : x_2});
    endrule

    rule rule_in_rsrel_00;
        $display ("Rule fired: rule_in_rsrel_00 at %t", $time);
        let x_0 <- getDLReady_00();
        let x_1 <- startRelease_00((x_0).r_id);
        Struct1 x_2 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        Struct6 x_3 = (Struct6 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_2,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id, ir_by_victim :
        Struct5 {valid : (Bool)'(False), data : unpack(0)}});
        let x_4 <- enq_fifoN2I_00(x_3);
    endrule

    rule rule_ir_cache_00;
        $display ("Rule fired: rule_ir_cache_00 at %t", $time);
        let x_0 <- deq_fifoN2I_00();
        when (! (((x_0).ir_by_victim).valid), noAction);
        Struct1 x_1 = ((x_0).ir_msg);
        let x_2 <- cache__00__infoRq((x_1).addr);
        let x_3 <- enq_fifoI2L_00(x_0);
    endrule

    rule rule_ir_victims_00;
        $display ("Rule fired: rule_ir_victims_00 at %t", $time);
        let x_0 <- deq_fifoN2I_00();
        when (((x_0).ir_by_victim).valid, noAction);
        let x_1 <- enq_fifoI2L_00(x_0);
    endrule

    rule rule_lr_cache_00;
        $display ("Rule fired: rule_lr_cache_00 at %t", $time);
        let x_0 <- deq_fifoI2L_00();
        when (! (((x_0).ir_by_victim).valid), noAction);
        let x_1 <- cache__00__infoRsValueRq(((x_0).ir_msg).addr);
        Struct12 x_2 = (Struct12 {lr_ir_pp : x_0, lr_ir : x_1, lr_value :
        unpack(0)});
        let x_3 <- enq_fifoL2E_00(x_2);
    endrule

    rule rule_lr_victims_00;
        $display ("Rule fired: rule_lr_victims_00 at %t", $time);
        let x_0 <- deq_fifoI2L_00();
        when (((x_0).ir_by_victim).valid, noAction);
        Bit#(3) x_1 = (((x_0).ir_by_victim).data);
        let x_2 <- victims__00__getVictim(x_1);
        Struct9 x_3 = (Struct9 {info_index : unpack(0), info_hit : unpack(0),
        info_way : unpack(0), edir_hit : unpack(0), edir_way : unpack(0),
        edir_slot : unpack(0), info : (x_2).victim_info, may_victim :
        unpack(0), reps : unpack(0)});
        Struct12 x_4 = (Struct12 {lr_ir_pp : x_0, lr_ir : x_3, lr_value :
        (x_2).victim_value});
        let x_5 <- enq_fifoL2E_00(x_4);
    endrule

    rule rule_exec_00_000000;
        $display ("Rule fired: rule_exec_00_000000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_14).dir_st))) && ((x_13) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))}).dir_excl)))},
        value_write : (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_20}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_001000;
        $display ("Rule fired: rule_exec_00_001000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) && (((x_14).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_01000;
        $display ("Rule fired: rule_exec_00_01000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_03000;
        $display ("Rule fired: rule_exec_00_03000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h8)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_10000;
        $display ("Rule fired: rule_exec_00_10000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) || (((x_13) ==
        ((Bit#(3))'(3'h2))) && (((x_12) == ((Bool)'(True))) &&
        ((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__00__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren00(x_23);
        let x_25 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_11000;
        $display ("Rule fired: rule_exec_00_11000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_14000;
        $display ("Rule fired: rule_exec_00_14000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h8)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_15000;
        $display ("Rule fired: rule_exec_00_15000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))) == ((Bit#(4))'(4'h0)))) && (((x_12) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_13))) &&
        (((x_14).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h8)});
        let x_20 <- broadcast_parentChildren00(Struct22 {cs_inds :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_25000;
        $display ("Rule fired: rule_exec_00_25000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2600000;
        $display ("Rule fired: rule_exec_00_2600000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2601000;
        $display ("Rule fired: rule_exec_00_2601000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_261000;
        $display ("Rule fired: rule_exec_00_261000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_27000;
        $display ("Rule fired: rule_exec_00_27000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_28000;
        $display ("Rule fired: rule_exec_00_28000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_290000;
        $display ("Rule fired: rule_exec_00_290000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_291000;
        $display ("Rule fired: rule_exec_00_291000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_210000;
        $display ("Rule fired: rule_exec_00_210000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_211000;
        $display ("Rule fired: rule_exec_00_211000 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        ((x_19).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_19).value_write, value :
        (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__00__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        Struct19 x_24 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_000001;
        $display ("Rule fired: rule_exec_00_000001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_14).dir_st))) && ((x_13) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))}).dir_excl)))},
        value_write : (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_20}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_001001;
        $display ("Rule fired: rule_exec_00_001001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) && (((x_14).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_01001;
        $display ("Rule fired: rule_exec_00_01001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_03001;
        $display ("Rule fired: rule_exec_00_03001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h9)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_10001;
        $display ("Rule fired: rule_exec_00_10001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) || (((x_13) ==
        ((Bit#(3))'(3'h2))) && (((x_12) == ((Bool)'(True))) &&
        ((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__00__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren00(x_23);
        let x_25 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_11001;
        $display ("Rule fired: rule_exec_00_11001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_14001;
        $display ("Rule fired: rule_exec_00_14001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h9)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_15001;
        $display ("Rule fired: rule_exec_00_15001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))) == ((Bit#(4))'(4'h0)))) && (((x_12) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_13))) &&
        (((x_14).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h9)});
        let x_20 <- broadcast_parentChildren00(Struct22 {cs_inds :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_25001;
        $display ("Rule fired: rule_exec_00_25001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2600001;
        $display ("Rule fired: rule_exec_00_2600001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2601001;
        $display ("Rule fired: rule_exec_00_2601001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_261001;
        $display ("Rule fired: rule_exec_00_261001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_27001;
        $display ("Rule fired: rule_exec_00_27001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_28001;
        $display ("Rule fired: rule_exec_00_28001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_290001;
        $display ("Rule fired: rule_exec_00_290001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_291001;
        $display ("Rule fired: rule_exec_00_291001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_210001;
        $display ("Rule fired: rule_exec_00_210001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_211001;
        $display ("Rule fired: rule_exec_00_211001 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        ((x_19).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_19).value_write, value :
        (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__00__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        Struct19 x_24 = (Struct19 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_000002;
        $display ("Rule fired: rule_exec_00_000002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_14).dir_st))) && ((x_13) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))}).dir_excl)))},
        value_write : (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_20}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_001002;
        $display ("Rule fired: rule_exec_00_001002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) && (((x_14).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_01002;
        $display ("Rule fired: rule_exec_00_01002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_03002;
        $display ("Rule fired: rule_exec_00_03002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'ha)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_10002;
        $display ("Rule fired: rule_exec_00_10002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) || (((x_13) ==
        ((Bit#(3))'(3'h2))) && (((x_12) == ((Bool)'(True))) &&
        ((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__00__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren00(x_23);
        let x_25 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_11002;
        $display ("Rule fired: rule_exec_00_11002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_14002;
        $display ("Rule fired: rule_exec_00_14002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'ha)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_15002;
        $display ("Rule fired: rule_exec_00_15002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))) == ((Bit#(4))'(4'h0)))) && (((x_12) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_13))) &&
        (((x_14).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'ha)});
        let x_20 <- broadcast_parentChildren00(Struct22 {cs_inds :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_25002;
        $display ("Rule fired: rule_exec_00_25002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2600002;
        $display ("Rule fired: rule_exec_00_2600002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2601002;
        $display ("Rule fired: rule_exec_00_2601002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_261002;
        $display ("Rule fired: rule_exec_00_261002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_27002;
        $display ("Rule fired: rule_exec_00_27002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_28002;
        $display ("Rule fired: rule_exec_00_28002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_290002;
        $display ("Rule fired: rule_exec_00_290002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_291002;
        $display ("Rule fired: rule_exec_00_291002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_210002;
        $display ("Rule fired: rule_exec_00_210002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_211002;
        $display ("Rule fired: rule_exec_00_211002 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        ((x_19).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_19).value_write, value :
        (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__00__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        Struct19 x_24 = (Struct19 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_000003;
        $display ("Rule fired: rule_exec_00_000003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_14).dir_st))) && ((x_13) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))}).dir_excl)))},
        value_write : (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_20}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_001003;
        $display ("Rule fired: rule_exec_00_001003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) && (((x_14).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_01003;
        $display ("Rule fired: rule_exec_00_01003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_03003;
        $display ("Rule fired: rule_exec_00_03003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'hb)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_10003;
        $display ("Rule fired: rule_exec_00_10003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) || (((x_13) ==
        ((Bit#(3))'(3'h2))) && (((x_12) == ((Bool)'(True))) &&
        ((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__00__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren00(x_23);
        let x_25 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_11003;
        $display ("Rule fired: rule_exec_00_11003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_13))) && (! (((Bit#(3))'(3'h2)) < ((x_14).dir_st)))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_00(Struct20 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_14003;
        $display ("Rule fired: rule_exec_00_14003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_13))) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'hb)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_15003;
        $display ("Rule fired: rule_exec_00_15003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))) == ((Bit#(4))'(4'h0)))) && (((x_12) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_13))) &&
        (((x_14).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'hb)});
        let x_20 <- broadcast_parentChildren00(Struct22 {cs_inds :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_25003;
        $display ("Rule fired: rule_exec_00_25003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2600003;
        $display ("Rule fired: rule_exec_00_2600003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_2601003;
        $display ("Rule fired: rule_exec_00_2601003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_261003;
        $display ("Rule fired: rule_exec_00_261003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_27003;
        $display ("Rule fired: rule_exec_00_27003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_28003;
        $display ("Rule fired: rule_exec_00_28003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_290003;
        $display ("Rule fired: rule_exec_00_290003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(False))) && (((((((x_14).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_14).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_291003;
        $display ("Rule fired: rule_exec_00_291003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_14).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_14).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_14).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_14).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (unpack(0))))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl,
        dir_sharers : ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__00__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_210003;
        $display ("Rule fired: rule_exec_00_210003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && (((x_13) == ((Bit#(3))'(3'h2)))
        && (((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) && (((x_14).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_14).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value, may_victim : (x_16).may_victim, reps :
        (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_211003;
        $display ("Rule fired: rule_exec_00_211003 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_14).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_14).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_14).dir_st) == ((Bit#(3))'(3'h3))) && (((x_14).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_14).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_14).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        ((x_19).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_19).value_write, value :
        (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__00__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        Struct19 x_24 = (Struct19 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_020;
        $display ("Rule fired: rule_exec_00_020 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct17 x_18 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_14).dir_excl, dir_sharers :
        (((x_14).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_14).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))}).dir_excl)))}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps : (x_19).reps});
        Struct17 x_21 = (Struct17 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_20).info).mesi_status, mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps : (x_20).reps});
        Struct17 x_22 = (Struct17 {addr : (x_21).addr, info_write :
        (x_21).info_write, info_hit : (x_21).info_hit, info_way :
        (x_21).info_way, edir_hit : (x_21).edir_hit, edir_way :
        (x_21).edir_way, edir_slot : (x_21).edir_slot, info : (x_21).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_21).may_victim, reps :
        (x_21).reps});
        let x_25 = ?;
        if ((x_8).valid) begin
            let x_23 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_22).info, victim_value :
            ((x_22).value_write ? ((x_22).value) : (x_9))});
            x_25 = x_9;
        end else begin
            let x_24 <- cache__00__valueRsLineRq(x_22);
            x_25 = x_24;
        end
        let x_26 <- releaseMSHR_00(x_4);
        Struct19 x_27 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_28 <- makeEnq_parentChildren00(x_27);
    endrule

    rule rule_exec_00_021;
        $display ("Rule fired: rule_exec_00_021 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct17 x_18 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_18).value_write, value :
        (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps : (x_19).reps});
        Struct17 x_21 = (Struct17 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_20).info).mesi_status, mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps : (x_20).reps});
        Struct17 x_22 = (Struct17 {addr : (x_21).addr, info_write :
        (x_21).info_write, info_hit : (x_21).info_hit, info_way :
        (x_21).info_way, edir_hit : (x_21).edir_hit, edir_way :
        (x_21).edir_way, edir_slot : (x_21).edir_slot, info : (x_21).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_21).may_victim, reps :
        (x_21).reps});
        let x_25 = ?;
        if ((x_8).valid) begin
            let x_23 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_22).info, victim_value :
            ((x_22).value_write ? ((x_22).value) : (x_9))});
            x_25 = x_9;
        end else begin
            let x_24 <- cache__00__valueRsLineRq(x_22);
            x_25 = x_24;
        end
        let x_26 <- releaseMSHR_00(x_4);
        Struct19 x_27 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_28 <- makeEnq_parentChildren00(x_27);
    endrule

    rule rule_exec_00_041;
        $display ("Rule fired: rule_exec_00_041 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((Bool)'(True), noAction);
        Struct23 x_15 = (Struct23 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_10).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_10).m_dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_10).m_dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_10).m_dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))))}, msg :
        ((x_10).m_dl_rss)[((((x_10).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_10).m_dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_10).m_dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_10).m_dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0)))))))))))))]});
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ((x_10).m_qidx);
        Struct17 x_18 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : ((unpack(0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st, mesi_dir_sharers : (((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        ((unpack(0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_st) ==
        ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : unpack(0), dir_sharers : ((unpack(0)) | (((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : ((unpack(0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_excl)))},
        value_write : (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps : (x_19).reps});
        Struct17 x_21 = (Struct17 {addr : (x_20).addr, info_write :
        (x_20).info_write, info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : (x_20).info,
        value_write : (Bool)'(True), value : ((x_15).msg).value, may_victim :
        (x_20).may_victim, reps : (x_20).reps});
        Struct17 x_22 = (Struct17 {addr : (x_21).addr, info_write :
        (Bool)'(True), info_hit : (x_21).info_hit, info_way :
        (x_21).info_way, edir_hit : (x_21).edir_hit, edir_way :
        (x_21).edir_way, edir_slot : (x_21).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_21).info).mesi_status,
        mesi_dir_st : ((x_21).info).mesi_dir_st, mesi_dir_sharers :
        ((x_21).info).mesi_dir_sharers}, value_write : (x_21).value_write,
        value : (x_21).value, may_victim : (x_21).may_victim, reps :
        (x_21).reps});
        let x_25 = ?;
        if ((x_8).valid) begin
            let x_23 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_22).info, victim_value :
            ((x_22).value_write ? ((x_22).value) : (x_9))});
            x_25 = x_9;
        end else begin
            let x_24 <- cache__00__valueRsLineRq(x_22);
            x_25 = x_24;
        end
        let x_26 <- releaseMSHR_00(x_4);
        Struct19 x_27 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_28 <- makeEnq_parentChildren00(x_27);
    endrule

    rule rule_exec_00_05;
        $display ("Rule fired: rule_exec_00_05 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_14).dir_st))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_06;
        $display ("Rule fired: rule_exec_00_06 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_13))) && ((!
        (((x_14).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_14).dir_st))))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h4)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_071;
        $display ("Rule fired: rule_exec_00_071 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((Bool)'(True), noAction);
        Struct23 x_15 = (Struct23 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_10).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_10).m_dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_10).m_dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_10).m_dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))))}, msg :
        ((x_10).m_dl_rss)[((((x_10).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_10).m_dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_10).m_dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_10).m_dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0)))))))))))))]});
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ((x_10).m_qidx);
        Struct17 x_18 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : (unpack(0)) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_st,
        mesi_dir_sharers : (((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        unpack(0), dir_sharers : (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct16 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps : (x_19).reps});
        Struct17 x_21 = (Struct17 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_20).info).mesi_status, mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps : (x_20).reps});
        Struct17 x_22 = (Struct17 {addr : (x_21).addr, info_write :
        (x_21).info_write, info_hit : (x_21).info_hit, info_way :
        (x_21).info_way, edir_hit : (x_21).edir_hit, edir_way :
        (x_21).edir_way, edir_slot : (x_21).edir_slot, info : (x_21).info,
        value_write : (Bool)'(True), value : ((x_15).msg).value, may_victim :
        (x_21).may_victim, reps :
        (x_21).reps});
        let x_25 = ?;
        if ((x_8).valid) begin
            let x_23 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_22).info, victim_value :
            ((x_22).value_write ? ((x_22).value) : (x_9))});
            x_25 = x_9;
        end else begin
            let x_24 <- cache__00__valueRsLineRq(x_22);
            x_25 = x_24;
        end
        let x_26 <- releaseMSHR_00(x_4);
        Struct19 x_27 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_28 <- makeEnq_parentChildren00(x_27);
    endrule

    rule rule_exec_00_12;
        $display ("Rule fired: rule_exec_00_12 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((((x_14).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_14).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_14).dir_sharers) == (((Bit#(4))'(4'h1))
        << (({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])})[1:0])))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct17 x_18 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_17)[1:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_18).value_write, value :
        (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : ((x_19).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps : (x_19).reps});
        Struct17 x_21 = (Struct17 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_20).info).mesi_status, mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps :
        (x_20).reps});
        let x_24 = ?;
        if ((x_8).valid) begin
            let x_22 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_21).info, victim_value :
            ((x_21).value_write ? ((x_21).value) : (x_9))});
            x_24 = x_9;
        end else begin
            let x_23 <- cache__00__valueRsLineRq(x_21);
            x_24 = x_23;
        end
        let x_25 <- releaseMSHR_00(x_4);
        Struct19 x_26 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_27 <- makeEnq_parentChildren00(x_26);
    endrule

    rule rule_exec_00_13;
        $display ("Rule fired: rule_exec_00_13 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])})[1:0])))) ==
        ((Bit#(4))'(4'h0)))) && (((x_14).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        Struct1 x_15 = ((x_10).m_msg);
        Bit#(4) x_16 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct17 x_17 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_17).info).mesi_status,
        mesi_dir_st : ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value, may_victim : (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        let x_22 <- transferUpDown_00(Struct24 {r_id : x_4, r_dl_rss_from :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((x_16)[1:0])))});
        let x_23 <- broadcast_parentChildren00(Struct22 {cs_inds :
        ((x_14).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((x_16)[1:0]))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_161;
        $display ("Rule fired: rule_exec_00_161 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = ((x_10).m_msg);
        Bit#(4) x_16 = ((x_10).m_qidx);
        Struct17 x_17 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value, may_victim : (x_17).may_victim, reps :
        (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_19).info).mesi_status, mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__00__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_00(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_26 <- makeEnq_parentChildren00(x_25);
    endrule

    rule rule_exec_00_170;
        $display ("Rule fired: rule_exec_00_170 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_14).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_171;
        $display ("Rule fired: rule_exec_00_171 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_13) < ((Bit#(3))'(3'h3)))) && (((x_14).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_17 = (Struct17 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__00__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_190;
        $display ("Rule fired: rule_exec_00_190 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_14).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (x_14).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_20 <- broadcast_parentChildren00(Struct22 {cs_inds :
        (x_14).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_191;
        $display ("Rule fired: rule_exec_00_191 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((x_14).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_14).dir_st)))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_14).dir_excl)})[1:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(4))'(4'h4)});
        Struct19 x_20 = (Struct19 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_14).dir_excl)})[1:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_192;
        $display ("Rule fired: rule_exec_00_192 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_14).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_15 = (x_3);
        Struct17 x_16 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__00__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerDL_00(Struct21 {r_id : x_4, r_dl_rss_from :
        (x_14).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_20 <- broadcast_parentChildren00(Struct22 {cs_inds :
        (x_14).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_11010;
        $display ("Rule fired: rule_exec_00_11010 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = ((x_10).m_msg);
        Bit#(4) x_16 = ((x_10).m_qidx);
        Struct17 x_17 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value, may_victim : (x_17).may_victim, reps :
        (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_19).info).mesi_status, mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__00__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_00(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_26 <- makeEnq_parentChildren00(x_25);
    endrule

    rule rule_exec_00_11011;
        $display ("Rule fired: rule_exec_00_11011 at %t", $time);
        let x_0 <- deq_fifoL2E_00();
        Struct6 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct5 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = ((x_10).m_msg);
        Bit#(4) x_16 = ((x_10).m_qidx);
        Struct17 x_17 = (Struct17 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct17 x_18 = (Struct17 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct16 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct16 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value, may_victim : (x_17).may_victim, reps :
        (x_17).reps});
        Struct17 x_19 = (Struct17 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct17 x_20 = (Struct17 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_19).info).mesi_status, mesi_dir_st : ((x_19).info).mesi_dir_st,
        mesi_dir_sharers : ((x_19).info).mesi_dir_sharers}, value_write :
        (x_19).value_write, value : (x_19).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__00__setVictim(Struct18 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__00__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_00(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_26 <- makeEnq_parentChildren00(x_25);
    endrule

    rule rule_exec_00_20;
        $display ("Rule fired: rule_exec_00_20 at %t", $time);
        let x_0 <- victims__00__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct15 x_5 = (Struct15 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_7) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_8))
        && ((x_8) < ((Bit#(3))'(3'h4)))) && (((x_9).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_11 <- makeEnq_parentChildren00(x_10);
        let x_12 <- setULImm_00(x_4);
        let x_13 <- victims__00__setVictimRq(Struct25 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    rule rule_exec_00_21;
        $display ("Rule fired: rule_exec_00_21 at %t", $time);
        let x_0 <- victims__00__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct15 x_5 = (Struct15 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when ((((x_9).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_7) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_8))) || (((x_7) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) && ((x_8) <
        ((Bit#(3))'(3'h3)))))), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_11 <- makeEnq_parentChildren00(x_10);
        let x_12 <- setULImm_00(x_4);
        let x_13 <- victims__00__setVictimRq(Struct25 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    rule rule_exec_00_23;
        $display ("Rule fired: rule_exec_00_23 at %t", $time);
        let x_0 <- victims__00__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct15 x_5 = (Struct15 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when ((((x_8) == ((Bit#(3))'(3'h1))) && (! (((x_9).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_8) == ((Bit#(3))'(3'h2))) && ((x_7) ==
        ((Bool)'(False)))), noAction);
        let x_10 <- canImm_00(x_1);
        let x_11 <- victims__00__releaseVictim(x_1);
    endrule

    // No methods in this module
endmodule

interface Module134;

endinterface

module mkModule134#(function Action victims__000__setVictimRq(Struct49 _),
    function ActionValue#(Bit#(3)) setULImm_000(Struct1 _),
    function ActionValue#(Struct44) victims__000__getFirstVictim(),
    function Action victims__000__setVictim(Struct48 _),
    function Action registerUL_000(Struct47 _),
    function Action makeEnq_parentChildren000(Struct19 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__000__valueRsLineRq(Struct46 _),
    function ActionValue#(Struct45) getMSHR_000(Bit#(3) _),
    function ActionValue#(Struct43) deq_fifoL2E_000(),
    function ActionValue#(Struct44) victims__000__getVictim(Bit#(2) _),
    function Action enq_fifoL2E_000(Struct43 _),
    function ActionValue#(Struct41) cache__000__infoRsValueRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoI2L_000(),
    function Action enq_fifoI2L_000(Struct40 _),
    function Action cache__000__infoRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoN2I_000(),
    function ActionValue#(Struct38) getCRqSlot_000(Struct37 _),
    function ActionValue#(Bool) victims__000__hasVictim(),
    function ActionValue#(Struct2) deq_fifoCRqInput_000(),
    function Action releaseMSHR_000(Bit#(3) _),
    function ActionValue#(Bit#(3)) victims__000__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct37) getWait_000(),
    function Action startRelease_000(Bit#(3) _),
    function ActionValue#(Bit#(3)) getULReady_000(Bit#(64) _),
    function Action enq_fifoN2I_000(Struct40 _),
    function ActionValue#(Struct39) victims__000__findVictim(Bit#(64) _),
    function ActionValue#(Struct38) getPRqSlot_000(Struct37 _),
    function ActionValue#(Struct2) deq_fifoPInput_000())
    (Module134);

    rule rule_in_prq_000;
        $display ("Rule fired: rule_in_prq_000 at %t", $time);
        let x_0 <- deq_fifoPInput_000();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_000(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).in_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- victims__000__findVictim((x_2).addr);
            Struct40 x_5 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id,
            ir_by_victim : x_4});
            let x_6 <- enq_fifoN2I_000(x_5);
        end else begin

        end
    endrule

    rule rule_in_prs_000;
        $display ("Rule fired: rule_in_prs_000 at %t", $time);
        let x_0 <- deq_fifoPInput_000();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- getULReady_000((x_2).addr);
        let x_4 <- startRelease_000(x_3);
        let x_5 <- victims__000__findVictim((x_2).addr);
        Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : x_3, ir_by_victim :
        x_5});
        let x_7 <- enq_fifoN2I_000(x_6);
    endrule

    rule rule_in_retry_000;
        $display ("Rule fired: rule_in_retry_000 at %t", $time);
        let x_0 <- getWait_000();
        Struct1 x_1 = ((x_0).r_msg);
        let x_2 <- victims__000__findVictim((x_1).addr);
        Struct40 x_3 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : (x_0).r_msg_from, ir_mshr_id : (x_0).r_id,
        ir_by_victim : x_2});
        let x_4 <- enq_fifoN2I_000(x_3);
    endrule

    rule rule_in_invrs_000;
        $display ("Rule fired: rule_in_invrs_000 at %t", $time);
        let x_0 <- deq_fifoPInput_000();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- getULReady_000((x_2).addr);
        let x_4 <- victims__000__releaseVictim((x_2).addr);
        let x_5 <- releaseMSHR_000(x_3);
    endrule

    rule rule_in_crq_000;
        $display ("Rule fired: rule_in_crq_000 at %t", $time);
        let x_0 <- deq_fifoCRqInput_000();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when (((x_1)[3:2]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- victims__000__hasVictim();
        when (! (x_3), noAction);
        let x_4 <- getCRqSlot_000(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_4).s_has_slot,
        noAction);
        if (! ((x_4).s_conflict)) begin
            let x_5 <- victims__000__findVictim((x_2).addr);
            Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_4).s_id,
            ir_by_victim : x_5});
            let x_7 <- enq_fifoN2I_000(x_6);
        end else begin

        end
    endrule

    rule rule_ir_cache_000;
        $display ("Rule fired: rule_ir_cache_000 at %t", $time);
        let x_0 <- deq_fifoN2I_000();
        when (! (((x_0).ir_by_victim).valid), noAction);
        Struct1 x_1 = ((x_0).ir_msg);
        let x_2 <- cache__000__infoRq((x_1).addr);
        let x_3 <- enq_fifoI2L_000(x_0);
    endrule

    rule rule_ir_victims_000;
        $display ("Rule fired: rule_ir_victims_000 at %t", $time);
        let x_0 <- deq_fifoN2I_000();
        when (((x_0).ir_by_victim).valid, noAction);
        let x_1 <- enq_fifoI2L_000(x_0);
    endrule

    rule rule_lr_cache_000;
        $display ("Rule fired: rule_lr_cache_000 at %t", $time);
        let x_0 <- deq_fifoI2L_000();
        when (! (((x_0).ir_by_victim).valid), noAction);
        let x_1 <- cache__000__infoRsValueRq(((x_0).ir_msg).addr);
        Struct43 x_2 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_1, lr_value :
        unpack(0)});
        let x_3 <- enq_fifoL2E_000(x_2);
    endrule

    rule rule_lr_victims_000;
        $display ("Rule fired: rule_lr_victims_000 at %t", $time);
        let x_0 <- deq_fifoI2L_000();
        when (((x_0).ir_by_victim).valid, noAction);
        Bit#(2) x_1 = (((x_0).ir_by_victim).data);
        let x_2 <- victims__000__getVictim(x_1);
        Struct41 x_3 = (Struct41 {info_index : unpack(0), info_hit :
        unpack(0), info_way : unpack(0), edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_2).victim_info,
        may_victim : unpack(0), reps : unpack(0)});
        Struct43 x_4 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_3, lr_value :
        (x_2).victim_value});
        let x_5 <- enq_fifoL2E_000(x_4);
    endrule

    rule rule_exec_000_00;
        $display ("Rule fired: rule_exec_000_00 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__000__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_18}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 <- releaseMSHR_000(x_4);
    endrule

    rule rule_exec_000_01;
        $display ("Rule fired: rule_exec_000_01 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__000__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_000(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
    endrule

    rule rule_exec_000_020;
        $display ("Rule fired: rule_exec_000_020 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__000__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_000(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren000(x_25);
    endrule

    rule rule_exec_000_021;
        $display ("Rule fired: rule_exec_000_021 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__000__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_000(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren000(x_25);
    endrule

    rule rule_exec_000_03;
        $display ("Rule fired: rule_exec_000_03 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__000__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 <- releaseMSHR_000(x_4);
    endrule

    rule rule_exec_000_100;
        $display ("Rule fired: rule_exec_000_100 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_13) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__000__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren000(x_23);
        let x_25 <- releaseMSHR_000(x_4);
    endrule

    rule rule_exec_000_101;
        $display ("Rule fired: rule_exec_000_101 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && ((x_13) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__000__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
        let x_23 <- releaseMSHR_000(x_4);
    endrule

    rule rule_exec_000_11;
        $display ("Rule fired: rule_exec_000_11 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__000__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_000(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
    endrule

    rule rule_exec_000_12;
        $display ("Rule fired: rule_exec_000_12 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (x_18).info_write, info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : (x_18).info,
        value_write : (Bool)'(True), value : (x_16).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_19).info).mesi_status,
        mesi_dir_st : ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        Struct46 x_21 = (Struct46 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : ((x_20).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps :
        (x_20).reps});
        let x_24 = ?;
        if ((x_8).valid) begin
            let x_22 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_21).info, victim_value :
            ((x_21).value_write ? ((x_21).value) : (x_9))});
            x_24 = x_9;
        end else begin
            let x_23 <- cache__000__valueRsLineRq(x_21);
            x_24 = x_23;
        end
        let x_25 <- releaseMSHR_000(x_4);
        Struct19 x_26 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_27 <- makeEnq_parentChildren000(x_26);
    endrule

    rule rule_exec_000_130;
        $display ("Rule fired: rule_exec_000_130 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__000__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 <- releaseMSHR_000(x_4);
    endrule

    rule rule_exec_000_131;
        $display ("Rule fired: rule_exec_000_131 at %t", $time);
        let x_0 <- deq_fifoL2E_000();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h8)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__000__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__000__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 <- releaseMSHR_000(x_4);
    endrule

    rule rule_exec_000_20;
        $display ("Rule fired: rule_exec_000_20 at %t", $time);
        let x_0 <- victims__000__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_11 <- makeEnq_parentChildren000(x_10);
        let x_12 <- setULImm_000(x_4);
        let x_13 <- victims__000__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    rule rule_exec_000_21;
        $display ("Rule fired: rule_exec_000_21 at %t", $time);
        let x_0 <- victims__000__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_11 <- makeEnq_parentChildren000(x_10);
        let x_12 <- setULImm_000(x_4);
        let x_13 <- victims__000__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    // No methods in this module
endmodule

interface Module135;

endinterface

module mkModule135#(function Action victims__001__setVictimRq(Struct49 _),
    function ActionValue#(Bit#(3)) setULImm_001(Struct1 _),
    function ActionValue#(Struct44) victims__001__getFirstVictim(),
    function Action victims__001__setVictim(Struct48 _),
    function Action registerUL_001(Struct47 _),
    function Action makeEnq_parentChildren001(Struct19 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__001__valueRsLineRq(Struct46 _),
    function ActionValue#(Struct45) getMSHR_001(Bit#(3) _),
    function ActionValue#(Struct43) deq_fifoL2E_001(),
    function ActionValue#(Struct44) victims__001__getVictim(Bit#(2) _),
    function Action enq_fifoL2E_001(Struct43 _),
    function ActionValue#(Struct41) cache__001__infoRsValueRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoI2L_001(),
    function Action enq_fifoI2L_001(Struct40 _),
    function Action cache__001__infoRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoN2I_001(),
    function ActionValue#(Struct38) getCRqSlot_001(Struct37 _),
    function ActionValue#(Bool) victims__001__hasVictim(),
    function ActionValue#(Struct2) deq_fifoCRqInput_001(),
    function Action releaseMSHR_001(Bit#(3) _),
    function ActionValue#(Bit#(3)) victims__001__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct37) getWait_001(),
    function Action startRelease_001(Bit#(3) _),
    function ActionValue#(Bit#(3)) getULReady_001(Bit#(64) _),
    function Action enq_fifoN2I_001(Struct40 _),
    function ActionValue#(Struct39) victims__001__findVictim(Bit#(64) _),
    function ActionValue#(Struct38) getPRqSlot_001(Struct37 _),
    function ActionValue#(Struct2) deq_fifoPInput_001())
    (Module135);

    rule rule_in_prq_001;
        $display ("Rule fired: rule_in_prq_001 at %t", $time);
        let x_0 <- deq_fifoPInput_001();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_001(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).in_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- victims__001__findVictim((x_2).addr);
            Struct40 x_5 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id,
            ir_by_victim : x_4});
            let x_6 <- enq_fifoN2I_001(x_5);
        end else begin

        end
    endrule

    rule rule_in_prs_001;
        $display ("Rule fired: rule_in_prs_001 at %t", $time);
        let x_0 <- deq_fifoPInput_001();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- getULReady_001((x_2).addr);
        let x_4 <- startRelease_001(x_3);
        let x_5 <- victims__001__findVictim((x_2).addr);
        Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : x_3, ir_by_victim :
        x_5});
        let x_7 <- enq_fifoN2I_001(x_6);
    endrule

    rule rule_in_retry_001;
        $display ("Rule fired: rule_in_retry_001 at %t", $time);
        let x_0 <- getWait_001();
        Struct1 x_1 = ((x_0).r_msg);
        let x_2 <- victims__001__findVictim((x_1).addr);
        Struct40 x_3 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : (x_0).r_msg_from, ir_mshr_id : (x_0).r_id,
        ir_by_victim : x_2});
        let x_4 <- enq_fifoN2I_001(x_3);
    endrule

    rule rule_in_invrs_001;
        $display ("Rule fired: rule_in_invrs_001 at %t", $time);
        let x_0 <- deq_fifoPInput_001();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- getULReady_001((x_2).addr);
        let x_4 <- victims__001__releaseVictim((x_2).addr);
        let x_5 <- releaseMSHR_001(x_3);
    endrule

    rule rule_in_crq_001;
        $display ("Rule fired: rule_in_crq_001 at %t", $time);
        let x_0 <- deq_fifoCRqInput_001();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when (((x_1)[3:2]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- victims__001__hasVictim();
        when (! (x_3), noAction);
        let x_4 <- getCRqSlot_001(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_4).s_has_slot,
        noAction);
        if (! ((x_4).s_conflict)) begin
            let x_5 <- victims__001__findVictim((x_2).addr);
            Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_4).s_id,
            ir_by_victim : x_5});
            let x_7 <- enq_fifoN2I_001(x_6);
        end else begin

        end
    endrule

    rule rule_ir_cache_001;
        $display ("Rule fired: rule_ir_cache_001 at %t", $time);
        let x_0 <- deq_fifoN2I_001();
        when (! (((x_0).ir_by_victim).valid), noAction);
        Struct1 x_1 = ((x_0).ir_msg);
        let x_2 <- cache__001__infoRq((x_1).addr);
        let x_3 <- enq_fifoI2L_001(x_0);
    endrule

    rule rule_ir_victims_001;
        $display ("Rule fired: rule_ir_victims_001 at %t", $time);
        let x_0 <- deq_fifoN2I_001();
        when (((x_0).ir_by_victim).valid, noAction);
        let x_1 <- enq_fifoI2L_001(x_0);
    endrule

    rule rule_lr_cache_001;
        $display ("Rule fired: rule_lr_cache_001 at %t", $time);
        let x_0 <- deq_fifoI2L_001();
        when (! (((x_0).ir_by_victim).valid), noAction);
        let x_1 <- cache__001__infoRsValueRq(((x_0).ir_msg).addr);
        Struct43 x_2 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_1, lr_value :
        unpack(0)});
        let x_3 <- enq_fifoL2E_001(x_2);
    endrule

    rule rule_lr_victims_001;
        $display ("Rule fired: rule_lr_victims_001 at %t", $time);
        let x_0 <- deq_fifoI2L_001();
        when (((x_0).ir_by_victim).valid, noAction);
        Bit#(2) x_1 = (((x_0).ir_by_victim).data);
        let x_2 <- victims__001__getVictim(x_1);
        Struct41 x_3 = (Struct41 {info_index : unpack(0), info_hit :
        unpack(0), info_way : unpack(0), edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_2).victim_info,
        may_victim : unpack(0), reps : unpack(0)});
        Struct43 x_4 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_3, lr_value :
        (x_2).victim_value});
        let x_5 <- enq_fifoL2E_001(x_4);
    endrule

    rule rule_exec_001_00;
        $display ("Rule fired: rule_exec_001_00 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__001__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_18}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 <- releaseMSHR_001(x_4);
    endrule

    rule rule_exec_001_01;
        $display ("Rule fired: rule_exec_001_01 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__001__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_001(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
    endrule

    rule rule_exec_001_020;
        $display ("Rule fired: rule_exec_001_020 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__001__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_001(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren001(x_25);
    endrule

    rule rule_exec_001_021;
        $display ("Rule fired: rule_exec_001_021 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__001__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_001(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren001(x_25);
    endrule

    rule rule_exec_001_03;
        $display ("Rule fired: rule_exec_001_03 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h9)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__001__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 <- releaseMSHR_001(x_4);
    endrule

    rule rule_exec_001_100;
        $display ("Rule fired: rule_exec_001_100 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_13) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__001__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren001(x_23);
        let x_25 <- releaseMSHR_001(x_4);
    endrule

    rule rule_exec_001_101;
        $display ("Rule fired: rule_exec_001_101 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && ((x_13) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__001__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
        let x_23 <- releaseMSHR_001(x_4);
    endrule

    rule rule_exec_001_11;
        $display ("Rule fired: rule_exec_001_11 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__001__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_001(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
    endrule

    rule rule_exec_001_12;
        $display ("Rule fired: rule_exec_001_12 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (x_18).info_write, info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : (x_18).info,
        value_write : (Bool)'(True), value : (x_16).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_19).info).mesi_status,
        mesi_dir_st : ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        Struct46 x_21 = (Struct46 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : ((x_20).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps :
        (x_20).reps});
        let x_24 = ?;
        if ((x_8).valid) begin
            let x_22 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_21).info, victim_value :
            ((x_21).value_write ? ((x_21).value) : (x_9))});
            x_24 = x_9;
        end else begin
            let x_23 <- cache__001__valueRsLineRq(x_21);
            x_24 = x_23;
        end
        let x_25 <- releaseMSHR_001(x_4);
        Struct19 x_26 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_27 <- makeEnq_parentChildren001(x_26);
    endrule

    rule rule_exec_001_130;
        $display ("Rule fired: rule_exec_001_130 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h9)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__001__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 <- releaseMSHR_001(x_4);
    endrule

    rule rule_exec_001_131;
        $display ("Rule fired: rule_exec_001_131 at %t", $time);
        let x_0 <- deq_fifoL2E_001();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h9)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__001__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__001__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 <- releaseMSHR_001(x_4);
    endrule

    rule rule_exec_001_20;
        $display ("Rule fired: rule_exec_001_20 at %t", $time);
        let x_0 <- victims__001__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_11 <- makeEnq_parentChildren001(x_10);
        let x_12 <- setULImm_001(x_4);
        let x_13 <- victims__001__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    rule rule_exec_001_21;
        $display ("Rule fired: rule_exec_001_21 at %t", $time);
        let x_0 <- victims__001__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_11 <- makeEnq_parentChildren001(x_10);
        let x_12 <- setULImm_001(x_4);
        let x_13 <- victims__001__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    // No methods in this module
endmodule

interface Module136;

endinterface

module mkModule136#(function Action victims__002__setVictimRq(Struct49 _),
    function ActionValue#(Bit#(3)) setULImm_002(Struct1 _),
    function ActionValue#(Struct44) victims__002__getFirstVictim(),
    function Action victims__002__setVictim(Struct48 _),
    function Action registerUL_002(Struct47 _),
    function Action makeEnq_parentChildren002(Struct19 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__002__valueRsLineRq(Struct46 _),
    function ActionValue#(Struct45) getMSHR_002(Bit#(3) _),
    function ActionValue#(Struct43) deq_fifoL2E_002(),
    function ActionValue#(Struct44) victims__002__getVictim(Bit#(2) _),
    function Action enq_fifoL2E_002(Struct43 _),
    function ActionValue#(Struct41) cache__002__infoRsValueRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoI2L_002(),
    function Action enq_fifoI2L_002(Struct40 _),
    function Action cache__002__infoRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoN2I_002(),
    function ActionValue#(Struct38) getCRqSlot_002(Struct37 _),
    function ActionValue#(Bool) victims__002__hasVictim(),
    function ActionValue#(Struct2) deq_fifoCRqInput_002(),
    function Action releaseMSHR_002(Bit#(3) _),
    function ActionValue#(Bit#(3)) victims__002__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct37) getWait_002(),
    function Action startRelease_002(Bit#(3) _),
    function ActionValue#(Bit#(3)) getULReady_002(Bit#(64) _),
    function Action enq_fifoN2I_002(Struct40 _),
    function ActionValue#(Struct39) victims__002__findVictim(Bit#(64) _),
    function ActionValue#(Struct38) getPRqSlot_002(Struct37 _),
    function ActionValue#(Struct2) deq_fifoPInput_002())
    (Module136);

    rule rule_in_prq_002;
        $display ("Rule fired: rule_in_prq_002 at %t", $time);
        let x_0 <- deq_fifoPInput_002();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h2))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_002(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).in_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- victims__002__findVictim((x_2).addr);
            Struct40 x_5 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id,
            ir_by_victim : x_4});
            let x_6 <- enq_fifoN2I_002(x_5);
        end else begin

        end
    endrule

    rule rule_in_prs_002;
        $display ("Rule fired: rule_in_prs_002 at %t", $time);
        let x_0 <- deq_fifoPInput_002();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h2))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- getULReady_002((x_2).addr);
        let x_4 <- startRelease_002(x_3);
        let x_5 <- victims__002__findVictim((x_2).addr);
        Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : x_3, ir_by_victim :
        x_5});
        let x_7 <- enq_fifoN2I_002(x_6);
    endrule

    rule rule_in_retry_002;
        $display ("Rule fired: rule_in_retry_002 at %t", $time);
        let x_0 <- getWait_002();
        Struct1 x_1 = ((x_0).r_msg);
        let x_2 <- victims__002__findVictim((x_1).addr);
        Struct40 x_3 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : (x_0).r_msg_from, ir_mshr_id : (x_0).r_id,
        ir_by_victim : x_2});
        let x_4 <- enq_fifoN2I_002(x_3);
    endrule

    rule rule_in_invrs_002;
        $display ("Rule fired: rule_in_invrs_002 at %t", $time);
        let x_0 <- deq_fifoPInput_002();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h2))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- getULReady_002((x_2).addr);
        let x_4 <- victims__002__releaseVictim((x_2).addr);
        let x_5 <- releaseMSHR_002(x_3);
    endrule

    rule rule_in_crq_002;
        $display ("Rule fired: rule_in_crq_002 at %t", $time);
        let x_0 <- deq_fifoCRqInput_002();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when (((x_1)[3:2]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- victims__002__hasVictim();
        when (! (x_3), noAction);
        let x_4 <- getCRqSlot_002(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_4).s_has_slot,
        noAction);
        if (! ((x_4).s_conflict)) begin
            let x_5 <- victims__002__findVictim((x_2).addr);
            Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_4).s_id,
            ir_by_victim : x_5});
            let x_7 <- enq_fifoN2I_002(x_6);
        end else begin

        end
    endrule

    rule rule_ir_cache_002;
        $display ("Rule fired: rule_ir_cache_002 at %t", $time);
        let x_0 <- deq_fifoN2I_002();
        when (! (((x_0).ir_by_victim).valid), noAction);
        Struct1 x_1 = ((x_0).ir_msg);
        let x_2 <- cache__002__infoRq((x_1).addr);
        let x_3 <- enq_fifoI2L_002(x_0);
    endrule

    rule rule_ir_victims_002;
        $display ("Rule fired: rule_ir_victims_002 at %t", $time);
        let x_0 <- deq_fifoN2I_002();
        when (((x_0).ir_by_victim).valid, noAction);
        let x_1 <- enq_fifoI2L_002(x_0);
    endrule

    rule rule_lr_cache_002;
        $display ("Rule fired: rule_lr_cache_002 at %t", $time);
        let x_0 <- deq_fifoI2L_002();
        when (! (((x_0).ir_by_victim).valid), noAction);
        let x_1 <- cache__002__infoRsValueRq(((x_0).ir_msg).addr);
        Struct43 x_2 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_1, lr_value :
        unpack(0)});
        let x_3 <- enq_fifoL2E_002(x_2);
    endrule

    rule rule_lr_victims_002;
        $display ("Rule fired: rule_lr_victims_002 at %t", $time);
        let x_0 <- deq_fifoI2L_002();
        when (((x_0).ir_by_victim).valid, noAction);
        Bit#(2) x_1 = (((x_0).ir_by_victim).data);
        let x_2 <- victims__002__getVictim(x_1);
        Struct41 x_3 = (Struct41 {info_index : unpack(0), info_hit :
        unpack(0), info_way : unpack(0), edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_2).victim_info,
        may_victim : unpack(0), reps : unpack(0)});
        Struct43 x_4 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_3, lr_value :
        (x_2).victim_value});
        let x_5 <- enq_fifoL2E_002(x_4);
    endrule

    rule rule_exec_002_00;
        $display ("Rule fired: rule_exec_002_00 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__002__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_18}});
        let x_20 <- makeEnq_parentChildren002(x_19);
        let x_21 <- releaseMSHR_002(x_4);
    endrule

    rule rule_exec_002_01;
        $display ("Rule fired: rule_exec_002_01 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__002__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_002(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren002(x_20);
    endrule

    rule rule_exec_002_020;
        $display ("Rule fired: rule_exec_002_020 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h2))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__002__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_002(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren002(x_25);
    endrule

    rule rule_exec_002_021;
        $display ("Rule fired: rule_exec_002_021 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h2))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__002__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_002(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren002(x_25);
    endrule

    rule rule_exec_002_03;
        $display ("Rule fired: rule_exec_002_03 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'ha)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__002__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren002(x_22);
        let x_24 <- releaseMSHR_002(x_4);
    endrule

    rule rule_exec_002_100;
        $display ("Rule fired: rule_exec_002_100 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_13) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__002__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren002(x_23);
        let x_25 <- releaseMSHR_002(x_4);
    endrule

    rule rule_exec_002_101;
        $display ("Rule fired: rule_exec_002_101 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && ((x_13) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__002__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren002(x_21);
        let x_23 <- releaseMSHR_002(x_4);
    endrule

    rule rule_exec_002_11;
        $display ("Rule fired: rule_exec_002_11 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__002__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_002(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren002(x_20);
    endrule

    rule rule_exec_002_12;
        $display ("Rule fired: rule_exec_002_12 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h2))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (x_18).info_write, info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : (x_18).info,
        value_write : (Bool)'(True), value : (x_16).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_19).info).mesi_status,
        mesi_dir_st : ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        Struct46 x_21 = (Struct46 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : ((x_20).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps :
        (x_20).reps});
        let x_24 = ?;
        if ((x_8).valid) begin
            let x_22 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_21).info, victim_value :
            ((x_21).value_write ? ((x_21).value) : (x_9))});
            x_24 = x_9;
        end else begin
            let x_23 <- cache__002__valueRsLineRq(x_21);
            x_24 = x_23;
        end
        let x_25 <- releaseMSHR_002(x_4);
        Struct19 x_26 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_27 <- makeEnq_parentChildren002(x_26);
    endrule

    rule rule_exec_002_130;
        $display ("Rule fired: rule_exec_002_130 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'ha)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__002__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren002(x_22);
        let x_24 <- releaseMSHR_002(x_4);
    endrule

    rule rule_exec_002_131;
        $display ("Rule fired: rule_exec_002_131 at %t", $time);
        let x_0 <- deq_fifoL2E_002();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_002(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'ha)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__002__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__002__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren002(x_22);
        let x_24 <- releaseMSHR_002(x_4);
    endrule

    rule rule_exec_002_20;
        $display ("Rule fired: rule_exec_002_20 at %t", $time);
        let x_0 <- victims__002__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_11 <- makeEnq_parentChildren002(x_10);
        let x_12 <- setULImm_002(x_4);
        let x_13 <- victims__002__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    rule rule_exec_002_21;
        $display ("Rule fired: rule_exec_002_21 at %t", $time);
        let x_0 <- victims__002__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_11 <- makeEnq_parentChildren002(x_10);
        let x_12 <- setULImm_002(x_4);
        let x_13 <- victims__002__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    // No methods in this module
endmodule

interface Module137;

endinterface

module mkModule137#(function Action victims__003__setVictimRq(Struct49 _),
    function ActionValue#(Bit#(3)) setULImm_003(Struct1 _),
    function ActionValue#(Struct44) victims__003__getFirstVictim(),
    function Action victims__003__setVictim(Struct48 _),
    function Action registerUL_003(Struct47 _),
    function Action makeEnq_parentChildren003(Struct19 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__003__valueRsLineRq(Struct46 _),
    function ActionValue#(Struct45) getMSHR_003(Bit#(3) _),
    function ActionValue#(Struct43) deq_fifoL2E_003(),
    function ActionValue#(Struct44) victims__003__getVictim(Bit#(2) _),
    function Action enq_fifoL2E_003(Struct43 _),
    function ActionValue#(Struct41) cache__003__infoRsValueRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoI2L_003(),
    function Action enq_fifoI2L_003(Struct40 _),
    function Action cache__003__infoRq(Bit#(64) _),
    function ActionValue#(Struct40) deq_fifoN2I_003(),
    function ActionValue#(Struct38) getCRqSlot_003(Struct37 _),
    function ActionValue#(Bool) victims__003__hasVictim(),
    function ActionValue#(Struct2) deq_fifoCRqInput_003(),
    function Action releaseMSHR_003(Bit#(3) _),
    function ActionValue#(Bit#(3)) victims__003__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct37) getWait_003(),
    function Action startRelease_003(Bit#(3) _),
    function ActionValue#(Bit#(3)) getULReady_003(Bit#(64) _),
    function Action enq_fifoN2I_003(Struct40 _),
    function ActionValue#(Struct39) victims__003__findVictim(Bit#(64) _),
    function ActionValue#(Struct38) getPRqSlot_003(Struct37 _),
    function ActionValue#(Struct2) deq_fifoPInput_003())
    (Module137);

    rule rule_in_prq_003;
        $display ("Rule fired: rule_in_prq_003 at %t", $time);
        let x_0 <- deq_fifoPInput_003();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h3))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_003(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).in_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- victims__003__findVictim((x_2).addr);
            Struct40 x_5 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id,
            ir_by_victim : x_4});
            let x_6 <- enq_fifoN2I_003(x_5);
        end else begin

        end
    endrule

    rule rule_in_prs_003;
        $display ("Rule fired: rule_in_prs_003 at %t", $time);
        let x_0 <- deq_fifoPInput_003();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h3))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- getULReady_003((x_2).addr);
        let x_4 <- startRelease_003(x_3);
        let x_5 <- victims__003__findVictim((x_2).addr);
        Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : x_3, ir_by_victim :
        x_5});
        let x_7 <- enq_fifoN2I_003(x_6);
    endrule

    rule rule_in_retry_003;
        $display ("Rule fired: rule_in_retry_003 at %t", $time);
        let x_0 <- getWait_003();
        Struct1 x_1 = ((x_0).r_msg);
        let x_2 <- victims__003__findVictim((x_1).addr);
        Struct40 x_3 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : (x_0).r_msg_from, ir_mshr_id : (x_0).r_id,
        ir_by_victim : x_2});
        let x_4 <- enq_fifoN2I_003(x_3);
    endrule

    rule rule_in_invrs_003;
        $display ("Rule fired: rule_in_invrs_003 at %t", $time);
        let x_0 <- deq_fifoPInput_003();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h3))}),
        noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- getULReady_003((x_2).addr);
        let x_4 <- victims__003__releaseVictim((x_2).addr);
        let x_5 <- releaseMSHR_003(x_3);
    endrule

    rule rule_in_crq_003;
        $display ("Rule fired: rule_in_crq_003 at %t", $time);
        let x_0 <- deq_fifoCRqInput_003();
        Bit#(4) x_1 = ((x_0).in_msg_from);
        when (((x_1)[3:2]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).in_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- victims__003__hasVictim();
        when (! (x_3), noAction);
        let x_4 <- getCRqSlot_003(Struct37 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_4).s_has_slot,
        noAction);
        if (! ((x_4).s_conflict)) begin
            let x_5 <- victims__003__findVictim((x_2).addr);
            Struct40 x_6 = (Struct40 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).in_msg, ir_msg_from : x_1, ir_mshr_id : (x_4).s_id,
            ir_by_victim : x_5});
            let x_7 <- enq_fifoN2I_003(x_6);
        end else begin

        end
    endrule

    rule rule_ir_cache_003;
        $display ("Rule fired: rule_ir_cache_003 at %t", $time);
        let x_0 <- deq_fifoN2I_003();
        when (! (((x_0).ir_by_victim).valid), noAction);
        Struct1 x_1 = ((x_0).ir_msg);
        let x_2 <- cache__003__infoRq((x_1).addr);
        let x_3 <- enq_fifoI2L_003(x_0);
    endrule

    rule rule_ir_victims_003;
        $display ("Rule fired: rule_ir_victims_003 at %t", $time);
        let x_0 <- deq_fifoN2I_003();
        when (((x_0).ir_by_victim).valid, noAction);
        let x_1 <- enq_fifoI2L_003(x_0);
    endrule

    rule rule_lr_cache_003;
        $display ("Rule fired: rule_lr_cache_003 at %t", $time);
        let x_0 <- deq_fifoI2L_003();
        when (! (((x_0).ir_by_victim).valid), noAction);
        let x_1 <- cache__003__infoRsValueRq(((x_0).ir_msg).addr);
        Struct43 x_2 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_1, lr_value :
        unpack(0)});
        let x_3 <- enq_fifoL2E_003(x_2);
    endrule

    rule rule_lr_victims_003;
        $display ("Rule fired: rule_lr_victims_003 at %t", $time);
        let x_0 <- deq_fifoI2L_003();
        when (((x_0).ir_by_victim).valid, noAction);
        Bit#(2) x_1 = (((x_0).ir_by_victim).data);
        let x_2 <- victims__003__getVictim(x_1);
        Struct41 x_3 = (Struct41 {info_index : unpack(0), info_hit :
        unpack(0), info_way : unpack(0), edir_hit : unpack(0), edir_way :
        unpack(0), edir_slot : unpack(0), info : (x_2).victim_info,
        may_victim : unpack(0), reps : unpack(0)});
        Struct43 x_4 = (Struct43 {lr_ir_pp : x_0, lr_ir : x_3, lr_value :
        (x_2).victim_value});
        let x_5 <- enq_fifoL2E_003(x_4);
    endrule

    rule rule_exec_003_00;
        $display ("Rule fired: rule_exec_003_00 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__003__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        Struct19 x_19 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_18}});
        let x_20 <- makeEnq_parentChildren003(x_19);
        let x_21 <- releaseMSHR_003(x_4);
    endrule

    rule rule_exec_003_01;
        $display ("Rule fired: rule_exec_003_01 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__003__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_003(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren003(x_20);
    endrule

    rule rule_exec_003_020;
        $display ("Rule fired: rule_exec_003_020 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h3))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__003__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_003(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren003(x_25);
    endrule

    rule rule_exec_003_021;
        $display ("Rule fired: rule_exec_003_021 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h3))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_19).may_victim, reps :
        (x_19).reps});
        let x_23 = ?;
        if ((x_8).valid) begin
            let x_21 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_20).info, victim_value :
            ((x_20).value_write ? ((x_20).value) : (x_9))});
            x_23 = x_9;
        end else begin
            let x_22 <- cache__003__valueRsLineRq(x_20);
            x_23 = x_22;
        end
        let x_24 <- releaseMSHR_003(x_4);
        Struct19 x_25 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (x_15).value}});
        let x_26 <- makeEnq_parentChildren003(x_25);
    endrule

    rule rule_exec_003_03;
        $display ("Rule fired: rule_exec_003_03 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'hb)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__003__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_21}});
        let x_23 <- makeEnq_parentChildren003(x_22);
        let x_24 <- releaseMSHR_003(x_4);
    endrule

    rule rule_exec_003_100;
        $display ("Rule fired: rule_exec_003_100 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_13) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps : (x_17).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_18).info).mesi_status,
        mesi_dir_st : ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value, may_victim : (x_18).may_victim, reps :
        (x_18).reps});
        let x_22 = ?;
        if ((x_8).valid) begin
            let x_20 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_19).info, victim_value :
            ((x_19).value_write ? ((x_19).value) : (x_9))});
            x_22 = x_9;
        end else begin
            let x_21 <- cache__003__valueRsLineRq(x_19);
            x_22 = x_21;
        end
        Struct19 x_23 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_24 <- makeEnq_parentChildren003(x_23);
        let x_25 <- releaseMSHR_003(x_4);
    endrule

    rule rule_exec_003_101;
        $display ("Rule fired: rule_exec_003_101 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12) == ((Bool)'(True))) && ((x_13) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_15).value, may_victim :
        (x_16).may_victim, reps :
        (x_16).reps});
        let x_20 = ?;
        if ((x_8).valid) begin
            let x_18 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_17).info, victim_value :
            ((x_17).value_write ? ((x_17).value) : (x_9))});
            x_20 = x_9;
        end else begin
            let x_19 <- cache__003__valueRsLineRq(x_17);
            x_20 = x_19;
        end
        Struct19 x_21 = (Struct19 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_22 <- makeEnq_parentChildren003(x_21);
        let x_23 <- releaseMSHR_003(x_4);
    endrule

    rule rule_exec_003_11;
        $display ("Rule fired: rule_exec_003_11 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_13)), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        let x_18 = ?;
        if ((x_8).valid) begin
            x_18 = x_9;
        end else begin
            let x_17 <- cache__003__valueRsLineRq(unpack(0));
            x_18 = x_17;
        end
        let x_19 <- registerUL_003(Struct47 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct19 x_20 = (Struct19 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren003(x_20);
    endrule

    rule rule_exec_003_12;
        $display ("Rule fired: rule_exec_003_12 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(2))'(2'h3))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((((x_10).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_10).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_10).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct1 x_16 = ((x_10).m_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),(((x_10).m_qidx)[1:0])});
        Struct46 x_18 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_19 = (Struct46 {addr : (x_18).addr, info_write :
        (x_18).info_write, info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : (x_18).info,
        value_write : (Bool)'(True), value : (x_16).value, may_victim :
        (x_18).may_victim, reps : (x_18).reps});
        Struct46 x_20 = (Struct46 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(True), mesi_status : ((x_19).info).mesi_status,
        mesi_dir_st : ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value, may_victim : (x_19).may_victim, reps :
        (x_19).reps});
        Struct46 x_21 = (Struct46 {addr : (x_20).addr, info_write :
        (Bool)'(True), info_hit : (x_20).info_hit, info_way :
        (x_20).info_way, edir_hit : (x_20).edir_hit, edir_way :
        (x_20).edir_way, edir_slot : (x_20).edir_slot, info : Struct10
        {mesi_owned : ((x_20).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_20).info).mesi_dir_st,
        mesi_dir_sharers : ((x_20).info).mesi_dir_sharers}, value_write :
        (x_20).value_write, value : (x_20).value, may_victim :
        (x_20).may_victim, reps :
        (x_20).reps});
        let x_24 = ?;
        if ((x_8).valid) begin
            let x_22 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_21).info, victim_value :
            ((x_21).value_write ? ((x_21).value) : (x_9))});
            x_24 = x_9;
        end else begin
            let x_23 <- cache__003__valueRsLineRq(x_21);
            x_24 = x_23;
        end
        let x_25 <- releaseMSHR_003(x_4);
        Struct19 x_26 = (Struct19 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_15).addr, value : unpack(0)}});
        let x_27 <- makeEnq_parentChildren003(x_26);
    endrule

    rule rule_exec_003_130;
        $display ("Rule fired: rule_exec_003_130 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'hb)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__003__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren003(x_22);
        let x_24 <- releaseMSHR_003(x_4);
    endrule

    rule rule_exec_003_131;
        $display ("Rule fired: rule_exec_003_131 at %t", $time);
        let x_0 <- deq_fifoL2E_003();
        Struct40 x_1 = ((x_0).lr_ir_pp);
        Bit#(4) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct41 x_6 = ((x_0).lr_ir);
        Struct10 x_7 = ((x_6).info);
        Struct39 x_8 = ((x_1).ir_by_victim);
        Vector#(4, Bit#(64)) x_9 = ((x_0).lr_value);
        let x_10 <- getMSHR_003(x_4);
        Vector#(4, Bit#(64)) x_11 = (unpack(0));
        Bool x_12 = ((x_7).mesi_owned);
        Bit#(3) x_13 = ((x_7).mesi_status);
        Struct16 x_14 = (Struct16 {dir_st : (((x_7).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_7).mesi_dir_st)),
        dir_excl : ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(4))'(4'hb)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_13) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_15 = (x_3);
        Struct46 x_16 = (Struct46 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0), may_victim : (x_6).may_victim, reps :
        (x_6).reps});
        Struct46 x_17 = (Struct46 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct10
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value, may_victim :
        (x_16).may_victim, reps : (x_16).reps});
        Struct46 x_18 = (Struct46 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct10
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value, may_victim :
        (x_17).may_victim, reps :
        (x_17).reps});
        let x_21 = ?;
        if ((x_8).valid) begin
            let x_19 <- victims__003__setVictim(Struct48 {victim_idx :
            (x_8).data, victim_info : (x_18).info, victim_value :
            ((x_18).value_write ? ((x_18).value) : (x_9))});
            x_21 = x_9;
        end else begin
            let x_20 <- cache__003__valueRsLineRq(x_18);
            x_21 = x_20;
        end
        Struct19 x_22 = (Struct19 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        unpack(0)}});
        let x_23 <- makeEnq_parentChildren003(x_22);
        let x_24 <- releaseMSHR_003(x_4);
    endrule

    rule rule_exec_003_20;
        $display ("Rule fired: rule_exec_003_20 at %t", $time);
        let x_0 <- victims__003__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_11 <- makeEnq_parentChildren003(x_10);
        let x_12 <- setULImm_003(x_4);
        let x_13 <- victims__003__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    rule rule_exec_003_21;
        $display ("Rule fired: rule_exec_003_21 at %t", $time);
        let x_0 <- victims__003__getFirstVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct10 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        Struct45 x_5 = (Struct45 {m_status : (Bit#(3))'(3'h5), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_6 = (unpack(0));
        Bool x_7 = ((x_2).mesi_owned);
        Bit#(3) x_8 = ((x_2).mesi_status);
        Struct16 x_9 = (Struct16 {dir_st : (((x_2).mesi_dir_st) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) : ((x_2).mesi_dir_st)),
        dir_excl : ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_2).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_2).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_2).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (unpack(0))))))))))))), dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        Struct19 x_10 = (Struct19 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_11 <- makeEnq_parentChildren003(x_10);
        let x_12 <- setULImm_003(x_4);
        let x_13 <- victims__003__setVictimRq(Struct49 {victim_addr : x_1,
        victim_req : x_12});
    endrule

    // No methods in this module
endmodule

// The CC interface is defined in the header part (thus in Header.bsv)

module mkCC#(function ActionValue#(Struct1) deq_fifo002(),
function Action enq_fifo001(Struct1 _),
function Action enq_fifo000(Struct1 _)) (CC);
    Module1 m1 <- mkModule1 ();
    Module2 m2 <- mkModule2 ();
    Module3 m3 <- mkModule3 ();
    Module4 m4 <- mkModule4 ();
    Module5 m5 <- mkModule5 ();
    Module6 m6 <- mkModule6 ();
    Module7 m7 <- mkModule7 ();
    Module8 m8 <- mkModule8 ();
    Module9 m9 <- mkModule9 ();
    Module10 m10 <- mkModule10 ();
    Module11 m11 <- mkModule11 ();
    Module12 m12 <- mkModule12 ();
    Module13 m13 <- mkModule13 ();
    Module14 m14 <- mkModule14 ();
    Module15 m15 <- mkModule15 ();
    Module16 m16 <- mkModule16 ();
    Module17 m17 <- mkModule17 ();
    Module18 m18 <- mkModule18 ();
    Module19 m19 <- mkModule19 ();
    Module20 m20 <- mkModule20 ();
    Module21 m21 <- mkModule21 ();
    Module22 m22 <- mkModule22 ();
    Module23 m23 <- mkModule23 ();
    Module24 m24 <- mkModule24 ();
    Module25 m25 <- mkModule25 ();
    Module26 m26 <- mkModule26 ();
    Module27 m27 <- mkModule27 ();
    Module28 m28 <- mkModule28 ();
    Module29 m29 <- mkModule29 ();
    Module30 m30 <- mkModule30 ();
    Module31 m31 <- mkModule31 ();
    Module32 m32 <- mkModule32 ();
    Module33 m33 <- mkModule33 ();
    Module34 m34 <- mkModule34 ();
    Module35 m35 <- mkModule35 ();
    Module36 m36 <- mkModule36 ();
    Module37 m37 <- mkModule37 ();
    Module38 m38 <- mkModule38 ();
    Module39 m39 <- mkModule39 ();
    Module40 m40 <- mkModule40 ();
    Module41 m41 <- mkModule41 ();
    Module42 m42 <- mkModule42 ();
    Module43 m43 <- mkModule43 ();
    Module44 m44 <- mkModule44 ();
    Module45 m45 <- mkModule45 ();
    Module46 m46 <- mkModule46 ();
    Module47 m47 <- mkModule47 ();
    Module48 m48 <- mkModule48 ();
    Module49 m49 <- mkModule49 ();
    Module50 m50 <- mkModule50 ();
    Module51 m51 <- mkModule51 ();
    Module52 m52 <- mkModule52 ();
    Module53 m53 <- mkModule53 ();
    Module54 m54 <- mkModule54 ();
    Module55 m55 <- mkModule55 ();
    Module56 m56 <- mkModule56 ();
    Module57 m57 <- mkModule57 ();
    Module58 m58 <- mkModule58 ();
    Module59 m59 <- mkModule59 ();
    Module60 m60 <- mkModule60 ();
    Module61 m61 <- mkModule61 ();
    Module62 m62 <- mkModule62 ();
    Module63 m63 <- mkModule63 ();
    Module64 m64 <- mkModule64 ();
    Module65 m65 <- mkModule65 ();
    Module66 m66 <- mkModule66 ();
    Module67 m67 <- mkModule67 ();
    Module68 m68 <- mkModule68 ();
    Module69 m69 <- mkModule69 ();
    Module70 m70 <- mkModule70 ();
    Module71 m71 <- mkModule71 ();
    Module72 m72 <- mkModule72 ();
    Module73 m73 <- mkModule73 ();
    Module74 m74 <- mkModule74 ();
    Module75 m75 <- mkModule75 ();
    Module76 m76 <- mkModule76 ();
    Module77 m77 <- mkModule77 ();
    Module78 m78 <- mkModule78 ();
    Module79 m79 <- mkModule79 ();
    Module80 m80 <- mkModule80 ();
    Module81 m81 <- mkModule81 ();
    Module82 m82 <- mkModule82 ();
    Module83 m83 <- mkModule83 ();
    Module84 m84 <- mkModule84 ();
    Module85 m85 <- mkModule85 ();
    Module86 m86 <- mkModule86 ();
    Module87 m87 <- mkModule87 ();
    Module88 m88 <- mkModule88 ();
    Module89 m89 <- mkModule89 ();
    Module90 m90 <- mkModule90 ();
    Module91 m91 <- mkModule91 ();
    Module92 m92 <- mkModule92 ();
    Module93 m93 <- mkModule93 ();
    Module94 m94 <- mkModule94 ();
    Module95 m95 <- mkModule95 ();
    Module96 m96 <- mkModule96 ();
    Module97 m97 <- mkModule97 ();
    Module98 m98 <- mkModule98 ();
    Module99 m99 <- mkModule99 ();
    Module100 m100 <- mkModule100 ();
    Module101 m101 <- mkModule101 ();
    Module102 m102 <- mkModule102 ();
    Module103 m103 <- mkModule103 ();
    Module104 m104 <- mkModule104 ();
    Module105 m105 <- mkModule105 ();
    Module106 m106 <- mkModule106 ();
    Module107 m107 <- mkModule107 (m94.deq_fifo0030, m76.deq_fifo0020,
    m58.deq_fifo0010, m1.enq_fifoCRqInput_00, m40.deq_fifo0000);
    Module108 m108 <- mkModule108 (m95.deq_fifo0031, m77.deq_fifo0021,
    m59.deq_fifo0011, m2.enq_fifoCRsInput_00, m41.deq_fifo0001);
    Module109 m109 <- mkModule109 (m3.enq_fifoPInput_00, deq_fifo002);

    Module110 m110 <- mkModule110 (m42.enq_fifo0002, m60.enq_fifo0012,
    m78.enq_fifo0022, m96.enq_fifo0032, enq_fifo001, enq_fifo000);
    Module111 m111 <- mkModule111 (m33.wrReq_repRam__00,
    m33.rdResp_repRam__00, m33.rdReq_repRam__00);
    Module112 m112 <- mkModule112 (m35.enq_fifoCRqInput_000,
    m43.deq_fifo00000);
    Module113 m113 <- mkModule113 (m36.enq_fifoPInput_000, m42.deq_fifo0002);

    Module114 m114 <- mkModule114 (m44.enq_fifo00002, m41.enq_fifo0001,
    m40.enq_fifo0000);
    Module115 m115 <- mkModule115 (m51.wrReq_repRam__000,
    m51.rdResp_repRam__000, m51.rdReq_repRam__000);
    Module116 m116 <- mkModule116 (m53.enq_fifoCRqInput_001,
    m61.deq_fifo00100);
    Module117 m117 <- mkModule117 (m54.enq_fifoPInput_001, m60.deq_fifo0012);

    Module118 m118 <- mkModule118 (m62.enq_fifo00102, m59.enq_fifo0011,
    m58.enq_fifo0010);
    Module119 m119 <- mkModule119 (m69.wrReq_repRam__001,
    m69.rdResp_repRam__001, m69.rdReq_repRam__001);
    Module120 m120 <- mkModule120 (m71.enq_fifoCRqInput_002,
    m79.deq_fifo00200);
    Module121 m121 <- mkModule121 (m72.enq_fifoPInput_002, m78.deq_fifo0022);

    Module122 m122 <- mkModule122 (m80.enq_fifo00202, m77.enq_fifo0021,
    m76.enq_fifo0020);
    Module123 m123 <- mkModule123 (m87.wrReq_repRam__002,
    m87.rdResp_repRam__002, m87.rdReq_repRam__002);
    Module124 m124 <- mkModule124 (m89.enq_fifoCRqInput_003,
    m97.deq_fifo00300);
    Module125 m125 <- mkModule125 (m90.enq_fifoPInput_003, m96.deq_fifo0032);

    Module126 m126 <- mkModule126 (m98.enq_fifo00302, m95.enq_fifo0031,
    m94.enq_fifo0030);
    Module127 m127 <- mkModule127 (m105.wrReq_repRam__003,
    m105.rdResp_repRam__003, m105.rdReq_repRam__003);
    Module128 m128 <- mkModule128 (m32.wrReq_dataRam__00,
    m24.wrReq_edirRam__00__7, m25.wrReq_edirRam__00__6,
    m26.wrReq_edirRam__00__5, m27.wrReq_edirRam__00__4,
    m28.wrReq_edirRam__00__3, m29.wrReq_edirRam__00__2,
    m30.wrReq_edirRam__00__1, m31.wrReq_edirRam__00__0, m111.repAccess__00,
    m7.victims__00__registerVictim, m8.wrReq_infoRam__00__15,
    m9.wrReq_infoRam__00__14, m10.wrReq_infoRam__00__13,
    m11.wrReq_infoRam__00__12, m12.wrReq_infoRam__00__11,
    m13.wrReq_infoRam__00__10, m14.wrReq_infoRam__00__9,
    m15.wrReq_infoRam__00__8, m16.wrReq_infoRam__00__7,
    m17.wrReq_infoRam__00__6, m18.wrReq_infoRam__00__5,
    m19.wrReq_infoRam__00__4, m20.wrReq_infoRam__00__3,
    m21.wrReq_infoRam__00__2, m22.wrReq_infoRam__00__1,
    m23.wrReq_infoRam__00__0, m32.rdResp_dataRam__00, m32.rdReq_dataRam__00,
    m111.repGetRs__00, m24.rdResp_edirRam__00__7, m25.rdResp_edirRam__00__6,
    m26.rdResp_edirRam__00__5, m27.rdResp_edirRam__00__4,
    m28.rdResp_edirRam__00__3, m29.rdResp_edirRam__00__2,
    m30.rdResp_edirRam__00__1, m31.rdResp_edirRam__00__0,
    m8.rdResp_infoRam__00__15, m9.rdResp_infoRam__00__14,
    m10.rdResp_infoRam__00__13, m11.rdResp_infoRam__00__12,
    m12.rdResp_infoRam__00__11, m13.rdResp_infoRam__00__10,
    m14.rdResp_infoRam__00__9, m15.rdResp_infoRam__00__8,
    m16.rdResp_infoRam__00__7, m17.rdResp_infoRam__00__6,
    m18.rdResp_infoRam__00__5, m19.rdResp_infoRam__00__4,
    m20.rdResp_infoRam__00__3, m21.rdResp_infoRam__00__2,
    m22.rdResp_infoRam__00__1, m23.rdResp_infoRam__00__0, m111.repGetRq__00,
    m24.rdReq_edirRam__00__7, m25.rdReq_edirRam__00__6,
    m26.rdReq_edirRam__00__5, m27.rdReq_edirRam__00__4,
    m28.rdReq_edirRam__00__3, m29.rdReq_edirRam__00__2,
    m30.rdReq_edirRam__00__1, m31.rdReq_edirRam__00__0,
    m8.rdReq_infoRam__00__15, m9.rdReq_infoRam__00__14,
    m10.rdReq_infoRam__00__13, m11.rdReq_infoRam__00__12,
    m12.rdReq_infoRam__00__11, m13.rdReq_infoRam__00__10,
    m14.rdReq_infoRam__00__9, m15.rdReq_infoRam__00__8,
    m16.rdReq_infoRam__00__7, m17.rdReq_infoRam__00__6,
    m18.rdReq_infoRam__00__5, m19.rdReq_infoRam__00__4,
    m20.rdReq_infoRam__00__3, m21.rdReq_infoRam__00__2,
    m22.rdReq_infoRam__00__1, m23.rdReq_infoRam__00__0);
    Module129 m129 <- mkModule129 (m50.wrReq_dataRam__000,
    m115.repAccess__000, m45.victims__000__registerVictim,
    m46.wrReq_infoRam__000__3, m47.wrReq_infoRam__000__2,
    m48.wrReq_infoRam__000__1, m49.wrReq_infoRam__000__0,
    m50.rdResp_dataRam__000, m50.rdReq_dataRam__000, m115.repGetRs__000,
    m46.rdResp_infoRam__000__3, m47.rdResp_infoRam__000__2,
    m48.rdResp_infoRam__000__1, m49.rdResp_infoRam__000__0,
    m115.repGetRq__000, m46.rdReq_infoRam__000__3, m47.rdReq_infoRam__000__2,
    m48.rdReq_infoRam__000__1, m49.rdReq_infoRam__000__0);
    Module130 m130 <- mkModule130 (m68.wrReq_dataRam__001,
    m119.repAccess__001, m63.victims__001__registerVictim,
    m64.wrReq_infoRam__001__3, m65.wrReq_infoRam__001__2,
    m66.wrReq_infoRam__001__1, m67.wrReq_infoRam__001__0,
    m68.rdResp_dataRam__001, m68.rdReq_dataRam__001, m119.repGetRs__001,
    m64.rdResp_infoRam__001__3, m65.rdResp_infoRam__001__2,
    m66.rdResp_infoRam__001__1, m67.rdResp_infoRam__001__0,
    m119.repGetRq__001, m64.rdReq_infoRam__001__3, m65.rdReq_infoRam__001__2,
    m66.rdReq_infoRam__001__1, m67.rdReq_infoRam__001__0);
    Module131 m131 <- mkModule131 (m86.wrReq_dataRam__002,
    m123.repAccess__002, m81.victims__002__registerVictim,
    m82.wrReq_infoRam__002__3, m83.wrReq_infoRam__002__2,
    m84.wrReq_infoRam__002__1, m85.wrReq_infoRam__002__0,
    m86.rdResp_dataRam__002, m86.rdReq_dataRam__002, m123.repGetRs__002,
    m82.rdResp_infoRam__002__3, m83.rdResp_infoRam__002__2,
    m84.rdResp_infoRam__002__1, m85.rdResp_infoRam__002__0,
    m123.repGetRq__002, m82.rdReq_infoRam__002__3, m83.rdReq_infoRam__002__2,
    m84.rdReq_infoRam__002__1, m85.rdReq_infoRam__002__0);
    Module132 m132 <- mkModule132 (m104.wrReq_dataRam__003,
    m127.repAccess__003, m99.victims__003__registerVictim,
    m100.wrReq_infoRam__003__3, m101.wrReq_infoRam__003__2,
    m102.wrReq_infoRam__003__1, m103.wrReq_infoRam__003__0,
    m104.rdResp_dataRam__003, m104.rdReq_dataRam__003, m127.repGetRs__003,
    m100.rdResp_infoRam__003__3, m101.rdResp_infoRam__003__2,
    m102.rdResp_infoRam__003__1, m103.rdResp_infoRam__003__0,
    m127.repGetRq__003, m100.rdReq_infoRam__003__3,
    m101.rdReq_infoRam__003__2, m102.rdReq_infoRam__003__1,
    m103.rdReq_infoRam__003__0);
    Module133 m133 <- mkModule133 (m34.canImm_00,
    m7.victims__00__setVictimRq, m34.setULImm_00,
    m7.victims__00__getFirstVictim, m34.transferUpDown_00,
    m110.broadcast_parentChildren00, m34.registerDL_00, m34.registerUL_00,
    m110.makeEnq_parentChildren00, m128.cache__00__valueRsLineRq,
    m7.victims__00__setVictim, m34.getMSHR_00, m6.deq_fifoL2E_00,
    m7.victims__00__getVictim, m6.enq_fifoL2E_00,
    m128.cache__00__infoRsValueRq, m5.deq_fifoI2L_00, m5.enq_fifoI2L_00,
    m128.cache__00__infoRq, m4.deq_fifoN2I_00, m34.getDLReady_00,
    m34.addRs_00, m2.deq_fifoCRsInput_00, m34.getCRqSlot_00,
    m7.victims__00__hasVictim, m1.deq_fifoCRqInput_00, m34.releaseMSHR_00,
    m7.victims__00__releaseVictim, m34.getWait_00, m34.startRelease_00,
    m34.getULReady_00, m4.enq_fifoN2I_00, m7.victims__00__findVictim,
    m34.getPRqSlot_00, m3.deq_fifoPInput_00);
    Module134 m134 <- mkModule134 (m45.victims__000__setVictimRq,
    m52.setULImm_000, m45.victims__000__getFirstVictim,
    m45.victims__000__setVictim, m52.registerUL_000,
    m114.makeEnq_parentChildren000, m129.cache__000__valueRsLineRq,
    m52.getMSHR_000, m39.deq_fifoL2E_000, m45.victims__000__getVictim,
    m39.enq_fifoL2E_000, m129.cache__000__infoRsValueRq, m38.deq_fifoI2L_000,
    m38.enq_fifoI2L_000, m129.cache__000__infoRq, m37.deq_fifoN2I_000,
    m52.getCRqSlot_000, m45.victims__000__hasVictim,
    m35.deq_fifoCRqInput_000, m52.releaseMSHR_000,
    m45.victims__000__releaseVictim, m52.getWait_000, m52.startRelease_000,
    m52.getULReady_000, m37.enq_fifoN2I_000, m45.victims__000__findVictim,
    m52.getPRqSlot_000, m36.deq_fifoPInput_000);
    Module135 m135 <- mkModule135 (m63.victims__001__setVictimRq,
    m70.setULImm_001, m63.victims__001__getFirstVictim,
    m63.victims__001__setVictim, m70.registerUL_001,
    m118.makeEnq_parentChildren001, m130.cache__001__valueRsLineRq,
    m70.getMSHR_001, m57.deq_fifoL2E_001, m63.victims__001__getVictim,
    m57.enq_fifoL2E_001, m130.cache__001__infoRsValueRq, m56.deq_fifoI2L_001,
    m56.enq_fifoI2L_001, m130.cache__001__infoRq, m55.deq_fifoN2I_001,
    m70.getCRqSlot_001, m63.victims__001__hasVictim,
    m53.deq_fifoCRqInput_001, m70.releaseMSHR_001,
    m63.victims__001__releaseVictim, m70.getWait_001, m70.startRelease_001,
    m70.getULReady_001, m55.enq_fifoN2I_001, m63.victims__001__findVictim,
    m70.getPRqSlot_001, m54.deq_fifoPInput_001);
    Module136 m136 <- mkModule136 (m81.victims__002__setVictimRq,
    m88.setULImm_002, m81.victims__002__getFirstVictim,
    m81.victims__002__setVictim, m88.registerUL_002,
    m122.makeEnq_parentChildren002, m131.cache__002__valueRsLineRq,
    m88.getMSHR_002, m75.deq_fifoL2E_002, m81.victims__002__getVictim,
    m75.enq_fifoL2E_002, m131.cache__002__infoRsValueRq, m74.deq_fifoI2L_002,
    m74.enq_fifoI2L_002, m131.cache__002__infoRq, m73.deq_fifoN2I_002,
    m88.getCRqSlot_002, m81.victims__002__hasVictim,
    m71.deq_fifoCRqInput_002, m88.releaseMSHR_002,
    m81.victims__002__releaseVictim, m88.getWait_002, m88.startRelease_002,
    m88.getULReady_002, m73.enq_fifoN2I_002, m81.victims__002__findVictim,
    m88.getPRqSlot_002, m72.deq_fifoPInput_002);
    Module137 m137 <- mkModule137 (m99.victims__003__setVictimRq,
    m106.setULImm_003, m99.victims__003__getFirstVictim,
    m99.victims__003__setVictim, m106.registerUL_003,
    m126.makeEnq_parentChildren003, m132.cache__003__valueRsLineRq,
    m106.getMSHR_003, m93.deq_fifoL2E_003, m99.victims__003__getVictim,
    m93.enq_fifoL2E_003, m132.cache__003__infoRsValueRq, m92.deq_fifoI2L_003,
    m92.enq_fifoI2L_003, m132.cache__003__infoRq, m91.deq_fifoN2I_003,
    m106.getCRqSlot_003, m99.victims__003__hasVictim,
    m89.deq_fifoCRqInput_003, m106.releaseMSHR_003,
    m99.victims__003__releaseVictim, m106.getWait_003, m106.startRelease_003,
    m106.getULReady_003, m91.enq_fifoN2I_003, m99.victims__003__findVictim,
    m106.getPRqSlot_003, m90.deq_fifoPInput_003);
    //// Interface

    function MemRqRs#(Struct1) getMemRqRs (function Action enq_rq (Struct1 _),
                                           function ActionValue#(Struct1) deq_rs ());
        return interface MemRqRs;
                   method mem_enq_rq = enq_rq;
                   method mem_deq_rs = deq_rs;
               endinterface;
    endfunction

    Vector#(L1Num, MemRqRs#(Struct1)) _l1Ifc = newVector();
    _l1Ifc[0] = getMemRqRs(m43.enq_fifo00000, m44.deq_fifo00002);
    _l1Ifc[1] = getMemRqRs(m61.enq_fifo00100, m62.deq_fifo00102);
    _l1Ifc[2] = getMemRqRs(m79.enq_fifo00200, m80.deq_fifo00202);
    _l1Ifc[3] = getMemRqRs(m97.enq_fifo00300, m98.deq_fifo00302);
    interface l1Ifc = _l1Ifc;

    interface DMA llDma;
        method dma_rdReq = m32.rdReq_dataRam__00;
        method dma_wrReq = m32.wrReq_dataRam__00;
        method dma_rdResp = m32.rdResp_dataRam__00;
    endinterface

endmodule
