CC_L1LL.bsv