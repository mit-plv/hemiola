CC_L1LL4.bsv