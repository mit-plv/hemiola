CCIfc2.bsv