import Vector::*;
import BuildVector::*;
import FIFO::*;
import FIFOF::*;
import RWBramCore::*;
import SpecialFIFOs::*;

typedef 4 L1Num;

interface MemRqRs;
    method Action mem_enq_rq (Struct1 rq);
    method ActionValue#(Struct1) mem_deq_rs ();
endinterface

interface DMA;
    method Action dma_rdReq (Bit#(14) addr);
    method Action dma_wrReq (Struct36 rq);
    method ActionValue#(Vector#(4, Bit#(64))) dma_rdResp ();
endinterface

interface CC;
    interface Vector#(L1Num, MemRqRs) l1Ifc;
    interface DMA llDma;
endinterface

typedef struct { Bit#(6) id; Bool type_; Bit#(64) addr; Vector#(4, Bit#(64)) value;  } Struct1 deriving(Eq, Bits);
typedef struct { Bool valid; Bit#(3) data;  } Struct10 deriving(Eq, Bits);
typedef struct { Bool mesi_owned; Bit#(3) mesi_status; Bit#(3) mesi_dir_st; Bit#(2) mesi_dir_sharers;  } Struct11 deriving(Eq, Bits);
typedef struct { Struct3 lr_ir_pp; Struct9 lr_ir;  } Struct12 deriving(Eq, Bits);
typedef struct { Bit#(2) m_status; Struct14 m_next; Bool m_is_ul; Struct1 m_msg; Bit#(3) m_qidx; Bool m_rsb; Bit#(2) m_dl_rss_from; Bit#(2) m_dl_rss_recv; Vector#(2, Struct1) m_dl_rss;  } Struct13 deriving(Eq, Bits);
typedef struct { Bool valid; Bit#(4) data;  } Struct14 deriving(Eq, Bits);
typedef struct { Bit#(3) dir_st; Bit#(1) dir_excl; Bit#(2) dir_sharers;  } Struct15 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_write; Bool info_hit; Bit#(4) info_way; Bool edir_hit; Bit#(3) edir_way; Struct10 edir_slot; Struct11 info; Bool value_write; Vector#(4, Bit#(64)) value;  } Struct16 deriving(Eq, Bits);
typedef struct { Bit#(2) enq_type; Bit#(1) enq_ch_idx; Struct1 enq_msg;  } Struct17 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bool r_ul_rsb; Bit#(1) r_ul_rsbTo;  } Struct18 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bit#(2) r_dl_rss_from; Bool r_dl_rsb; Bit#(3) r_dl_rsbTo;  } Struct19 deriving(Eq, Bits);
typedef struct { Bit#(1) ch_idx; Struct1 ch_msg;  } Struct2 deriving(Eq, Bits);
typedef struct { Bit#(2) cs_inds; Struct1 cs_msg;  } Struct20 deriving(Eq, Bits);
typedef struct { Bit#(3) cidx; Struct1 msg;  } Struct21 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bit#(2) r_dl_rss_from;  } Struct22 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(64) victim_addr; Struct11 victim_info; Vector#(4, Bit#(64)) victim_value; Struct14 victim_req;  } Struct23 deriving(Eq, Bits);
typedef struct { Bit#(64) victim_addr; Bit#(4) victim_req;  } Struct24 deriving(Eq, Bits);
typedef struct { Bit#(49) tag; Bit#(10) index; Struct26 victim_found;  } Struct25 deriving(Eq, Bits);
typedef struct { Bool valid; Bit#(1) data;  } Struct26 deriving(Eq, Bits);
typedef struct { Struct26 victim_found; Struct28 may_victim; Vector#(16, Bit#(8)) reps;  } Struct27 deriving(Eq, Bits);
typedef struct { Bit#(64) mv_addr; Struct11 mv_info;  } Struct28 deriving(Eq, Bits);
typedef struct { Bit#(49) tag; Struct11 value;  } Struct29 deriving(Eq, Bits);
typedef struct { Bool ir_is_rs_rel; Struct1 ir_msg; Bit#(3) ir_msg_from; Bit#(4) ir_mshr_id;  } Struct3 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(4) tm_way; Struct11 tm_value;  } Struct30 deriving(Eq, Bits);
typedef struct { Bit#(49) tag; Struct32 value;  } Struct31 deriving(Eq, Bits);
typedef struct { Bit#(3) mesi_edir_st; Bit#(2) mesi_edir_sharers;  } Struct32 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(3) tm_way; Struct32 tm_value;  } Struct33 deriving(Eq, Bits);
typedef struct { Bit#(10) addr; Struct29 datain;  } Struct34 deriving(Eq, Bits);
typedef struct { Bit#(1) acc_type; Vector#(16, Bit#(8)) acc_reps; Bit#(10) acc_index; Bit#(4) acc_way;  } Struct35 deriving(Eq, Bits);
typedef struct { Bit#(14) addr; Vector#(4, Bit#(64)) datain;  } Struct36 deriving(Eq, Bits);
typedef struct { Bit#(10) addr; Struct31 datain;  } Struct37 deriving(Eq, Bits);
typedef struct { Bool valid; Struct23 data;  } Struct38 deriving(Eq, Bits);
typedef struct { Bit#(10) addr; Vector#(16, Bit#(8)) datain;  } Struct39 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Struct1 r_msg; Bit#(3) r_msg_from;  } Struct4 deriving(Eq, Bits);
typedef struct { Bit#(9) info_index; Bool info_hit; Bit#(3) info_way; Bool edir_hit; Bit#(2) edir_way; Struct41 edir_slot; Struct11 info;  } Struct40 deriving(Eq, Bits);
typedef struct { Bool valid; Bit#(2) data;  } Struct41 deriving(Eq, Bits);
typedef struct { Struct3 lr_ir_pp; Struct40 lr_ir;  } Struct42 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_write; Bool info_hit; Bit#(3) info_way; Bool edir_hit; Bit#(2) edir_way; Struct41 edir_slot; Struct11 info; Bool value_write; Vector#(4, Bit#(64)) value;  } Struct43 deriving(Eq, Bits);
typedef struct { Bit#(50) tag; Bit#(9) index; Struct26 victim_found;  } Struct44 deriving(Eq, Bits);
typedef struct { Struct26 victim_found; Struct28 may_victim; Vector#(8, Bit#(8)) reps;  } Struct45 deriving(Eq, Bits);
typedef struct { Bit#(50) tag; Struct11 value;  } Struct46 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(3) tm_way; Struct11 tm_value;  } Struct47 deriving(Eq, Bits);
typedef struct { Bit#(50) tag; Struct32 value;  } Struct48 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(2) tm_way; Struct32 tm_value;  } Struct49 deriving(Eq, Bits);
typedef struct { Bool s_has_slot; Bool s_conflict; Bit#(4) s_id;  } Struct5 deriving(Eq, Bits);
typedef struct { Bit#(9) addr; Struct46 datain;  } Struct50 deriving(Eq, Bits);
typedef struct { Bit#(1) acc_type; Vector#(8, Bit#(8)) acc_reps; Bit#(9) acc_index; Bit#(3) acc_way;  } Struct51 deriving(Eq, Bits);
typedef struct { Bit#(12) addr; Vector#(4, Bit#(64)) datain;  } Struct52 deriving(Eq, Bits);
typedef struct { Bit#(9) addr; Struct48 datain;  } Struct53 deriving(Eq, Bits);
typedef struct { Bit#(9) addr; Vector#(8, Bit#(8)) datain;  } Struct54 deriving(Eq, Bits);
typedef struct { Bool ir_is_rs_rel; Struct1 ir_msg; Bit#(3) ir_msg_from; Bit#(3) ir_mshr_id;  } Struct55 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Struct1 r_msg; Bit#(3) r_msg_from;  } Struct56 deriving(Eq, Bits);
typedef struct { Bool s_has_slot; Bool s_conflict; Bit#(3) s_id;  } Struct57 deriving(Eq, Bits);
typedef struct { Bool valid; Struct56 data;  } Struct58 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bit#(64) r_addr;  } Struct59 deriving(Eq, Bits);
typedef struct { Bit#(1) r_dl_midx; Struct1 r_dl_msg;  } Struct6 deriving(Eq, Bits);
typedef struct { Bit#(8) info_index; Bool info_hit; Bit#(2) info_way; Bool edir_hit; void edir_way; Struct61 edir_slot; Struct11 info;  } Struct60 deriving(Eq, Bits);
typedef struct { Bool valid; void data;  } Struct61 deriving(Eq, Bits);
typedef struct { Struct55 lr_ir_pp; Struct60 lr_ir;  } Struct62 deriving(Eq, Bits);
typedef struct { Bit#(2) m_status; Struct10 m_next; Bool m_is_ul; Struct1 m_msg; Bit#(3) m_qidx; Bool m_rsb; Bit#(2) m_dl_rss_from; Bit#(2) m_dl_rss_recv; Vector#(2, Struct1) m_dl_rss;  } Struct63 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_write; Bool info_hit; Bit#(2) info_way; Bool edir_hit; void edir_way; Struct61 edir_slot; Struct11 info; Bool value_write; Vector#(4, Bit#(64)) value;  } Struct64 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bool r_ul_rsb; Bit#(1) r_ul_rsbTo;  } Struct65 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(64) victim_addr; Struct11 victim_info; Vector#(4, Bit#(64)) victim_value; Struct10 victim_req;  } Struct66 deriving(Eq, Bits);
typedef struct { Bit#(64) victim_addr; Bit#(3) victim_req;  } Struct67 deriving(Eq, Bits);
typedef struct { Bit#(51) tag; Bit#(8) index; Struct26 victim_found;  } Struct68 deriving(Eq, Bits);
typedef struct { Struct26 victim_found; Struct28 may_victim; Vector#(4, Bit#(8)) reps;  } Struct69 deriving(Eq, Bits);
typedef struct { Bool valid; Struct4 data;  } Struct7 deriving(Eq, Bits);
typedef struct { Bit#(51) tag; Struct11 value;  } Struct70 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(2) tm_way; Struct11 tm_value;  } Struct71 deriving(Eq, Bits);
typedef struct { Bit#(8) addr; Struct70 datain;  } Struct72 deriving(Eq, Bits);
typedef struct { Bit#(10) addr; Vector#(4, Bit#(64)) datain;  } Struct73 deriving(Eq, Bits);
typedef struct { Bit#(1) acc_type; Vector#(4, Bit#(8)) acc_reps; Bit#(8) acc_index; Bit#(2) acc_way;  } Struct74 deriving(Eq, Bits);
typedef struct { Bool valid; Struct66 data;  } Struct75 deriving(Eq, Bits);
typedef struct { Bit#(8) addr; Vector#(4, Bit#(8)) datain;  } Struct76 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bit#(2) r_dl_rss_from; Bool r_dl_rsb; Bit#(3) r_dl_rsbTo;  } Struct77 deriving(Eq, Bits);
typedef struct { Bit#(3) r_id; Bit#(2) r_dl_rss_from;  } Struct78 deriving(Eq, Bits);
typedef struct { Bit#(4) r_id; Bit#(64) r_addr;  } Struct8 deriving(Eq, Bits);
typedef struct { Bit#(10) info_index; Bool info_hit; Bit#(4) info_way; Bool edir_hit; Bit#(3) edir_way; Struct10 edir_slot; Struct11 info;  } Struct9 deriving(Eq, Bits);

interface Module1;
    method Action enq_fifoCRqInput00 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput00 ();
endinterface

module mkModule1 (Module1);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifoCRqInput00 (Struct2 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput00 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module2;
    method Action enq_fifoCRsInput00 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRsInput00 ();
endinterface

module mkModule2 (Module2);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifoCRsInput00 (Struct2 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifoCRsInput00 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module3;
    method Action enq_fifoInput00 (Struct3 x_0);
    method ActionValue#(Struct3) deq_fifoInput00 ();
endinterface

module mkModule3 (Module3);
    FIFOF#(Struct3) pff <- mkFIFOF();

    method Action enq_fifoInput00 (Struct3 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct3) deq_fifoInput00 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module4;
    method Action enq_fifoI2L00 (Struct3 x_0);
    method ActionValue#(Struct3) deq_fifoI2L00 ();
endinterface

module mkModule4 (Module4);
    FIFOF#(Struct3) pff <- mkFIFOF();

    method Action enq_fifoI2L00 (Struct3 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct3) deq_fifoI2L00 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module5;
    method Action enq_fifoL2E00 (Struct12 x_0);
    method ActionValue#(Struct12) deq_fifoL2E00 ();
endinterface

module mkModule5 (Module5);
    FIFOF#(Struct12) pff <- mkFIFOF();

    method Action enq_fifoL2E00 (Struct12 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct12) deq_fifoL2E00 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module6;
    method Action enq_cp_1__00 (Struct25 x_0);
    method ActionValue#(Struct25) deq_cp_1__00 ();
endinterface

module mkModule6 (Module6);
    FIFOF#(Struct25) pff <- mkPipelineFIFOF();

    method Action enq_cp_1__00 (Struct25 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct25) deq_cp_1__00 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module7;
    method Action enq_cp_2__00 (Struct27 x_0);
    method ActionValue#(Struct27) deq_cp_2__00 ();
endinterface

module mkModule7 (Module7);
    FIFOF#(Struct27) pff <- mkPipelineFIFOF();

    method Action enq_cp_2__00 (Struct27 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct27) deq_cp_2__00 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module8;
    method Action rdReq_infoRam__00__15 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__15 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__15 ();
endinterface

module mkModule8 (Module8);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'hf, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__15 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__15 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__15 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module9;
    method Action rdReq_infoRam__00__14 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__14 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__14 ();
endinterface

module mkModule9 (Module9);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'he, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__14 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__14 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__14 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module10;
    method Action rdReq_infoRam__00__13 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__13 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__13 ();
endinterface

module mkModule10 (Module10);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'hd, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__13 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__13 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__13 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module11;
    method Action rdReq_infoRam__00__12 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__12 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__12 ();
endinterface

module mkModule11 (Module11);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'hc, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__12 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__12 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__12 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module12;
    method Action rdReq_infoRam__00__11 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__11 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__11 ();
endinterface

module mkModule12 (Module12);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'hb, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__11 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__11 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__11 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module13;
    method Action rdReq_infoRam__00__10 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__10 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__10 ();
endinterface

module mkModule13 (Module13);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'ha, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__10 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__10 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__10 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module14;
    method Action rdReq_infoRam__00__9 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__9 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__9 ();
endinterface

module mkModule14 (Module14);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h9, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__9 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__9 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__9 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module15;
    method Action rdReq_infoRam__00__8 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__8 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__8 ();
endinterface

module mkModule15 (Module15);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h8, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__8 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__8 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__8 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module16;
    method Action rdReq_infoRam__00__7 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__7 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__7 ();
endinterface

module mkModule16 (Module16);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h7, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__7 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__7 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__7 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module17;
    method Action rdReq_infoRam__00__6 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__6 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__6 ();
endinterface

module mkModule17 (Module17);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h6, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__6 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__6 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__6 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module18;
    method Action rdReq_infoRam__00__5 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__5 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__5 ();
endinterface

module mkModule18 (Module18);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h5, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__5 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__5 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__5 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module19;
    method Action rdReq_infoRam__00__4 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__4 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__4 ();
endinterface

module mkModule19 (Module19);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h4, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__4 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__4 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__4 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module20;
    method Action rdReq_infoRam__00__3 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__3 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__3 ();
endinterface

module mkModule20 (Module20);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h3, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__3 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__3 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module21;
    method Action rdReq_infoRam__00__2 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__2 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__2 ();
endinterface

module mkModule21 (Module21);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h2, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__2 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__2 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module22;
    method Action rdReq_infoRam__00__1 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__1 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__1 ();
endinterface

module mkModule22 (Module22);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h1, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__1 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__1 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module23;
    method Action rdReq_infoRam__00__0 (Bit#(10) x_0);
    method Action wrReq_infoRam__00__0 (Struct34 x_0);
    method ActionValue#(Struct29) rdResp_infoRam__00__0 ();
endinterface

module mkModule23 (Module23);
    RWBramCore#(Bit#(10), Struct29) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct29 {tag: 49'h0, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__00__0 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__00__0 (Struct34 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct29) rdResp_infoRam__00__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module24;
    method Action rdReq_edirRam__00__7 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__7 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__7 ();
endinterface

module mkModule24 (Module24);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h7, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__7 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__7 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__7 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module25;
    method Action rdReq_edirRam__00__6 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__6 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__6 ();
endinterface

module mkModule25 (Module25);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h6, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__6 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__6 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__6 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module26;
    method Action rdReq_edirRam__00__5 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__5 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__5 ();
endinterface

module mkModule26 (Module26);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h5, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__5 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__5 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__5 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module27;
    method Action rdReq_edirRam__00__4 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__4 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__4 ();
endinterface

module mkModule27 (Module27);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h4, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__4 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__4 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__4 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module28;
    method Action rdReq_edirRam__00__3 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__3 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__3 ();
endinterface

module mkModule28 (Module28);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h3, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__3 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__3 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module29;
    method Action rdReq_edirRam__00__2 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__2 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__2 ();
endinterface

module mkModule29 (Module29);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h2, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__2 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__2 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module30;
    method Action rdReq_edirRam__00__1 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__1 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__1 ();
endinterface

module mkModule30 (Module30);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h1, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__1 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__1 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module31;
    method Action rdReq_edirRam__00__0 (Bit#(10) x_0);
    method Action wrReq_edirRam__00__0 (Struct37 x_0);
    method ActionValue#(Struct31) rdResp_edirRam__00__0 ();
endinterface

module mkModule31 (Module31);
    RWBramCore#(Bit#(10), Struct31) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct31 {tag: 49'h0, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__00__0 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__00__0 (Struct37 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct31) rdResp_edirRam__00__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module32;
    method Action rdReq_dataRam__00 (Bit#(14) x_0);
    method Action wrReq_dataRam__00 (Struct36 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__00 ();
endinterface

module mkModule32 (Module32);
    RWBramCore#(Bit#(14), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(14)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__00 (Bit#(14) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__00 (Struct36 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__00 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module33;
    method Action rdReq_repRam__00 (Bit#(10) x_0);
    method Action wrReq_repRam__00 (Struct39 x_0);
    method ActionValue#(Vector#(16, Bit#(8))) rdResp_repRam__00 ();
endinterface

module mkModule33 (Module33);
    RWBramCore#(Bit#(10), Vector#(16, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__00 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__00 (Struct39 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(16, Bit#(8))) rdResp_repRam__00 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module34;
    method ActionValue#(Struct13) getMSHR_00 (Bit#(4) x_0);
    method ActionValue#(Struct5) getPRqSlot_00 (Struct4 x_0);
    method ActionValue#(Struct5) getCRqSlot_00 (Struct4 x_0);
    method ActionValue#(Struct7) getWait_00 ();
    method Action registerUL_00 (Struct18 x_0);
    method Action registerDL_00 (Struct19 x_0);
    method ActionValue#(Bit#(4)) getULImm_00 (Struct1 x_0);
    method ActionValue#(Bit#(4)) getULCount_00 ();
    method Action transferUpDown_00 (Struct22 x_0);
    method ActionValue#(Bit#(4)) findUL_00 (Bit#(64) x_0);
    method ActionValue#(Bit#(4)) findDL_00 (Bit#(64) x_0);
    method Action releaseMSHR_00 (Bit#(4) x_0);
    method Action addRs_00 (Struct6 x_0);
    method ActionValue#(Struct8) getRsReady_00 ();
endinterface

module mkModule34
    (Module34);
    Reg#(Vector#(16, Struct13)) rqs_00 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct13) getMSHR_00 (Bit#(4) x_0);
        let x_1 = (rqs_00);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct5) getPRqSlot_00 (Struct4 x_0);
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (((((x_1)[(Bit#(4))'(4'hc)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hc)}) : (((((x_1)[(Bit#(4))'(4'hd)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hd)}) : (((((x_1)[(Bit#(4))'(4'he)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'he)}) : (((((x_1)[(Bit#(4))'(4'hf)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hf)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))))))))))))))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct14 x_6 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hc)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hc)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hc)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hc)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hd)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hd)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hd)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hd)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'he)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'he)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'he)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'he)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hf)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hf)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hf)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hf)}) : (Struct14 {valid
        : (Bool)'(False), data :
        unpack(0)})))))))))))))))))))))))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(4) x_8 = ((x_6).data);
        Struct5 x_9 = (Struct5 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct13 x_10 = ((x_1)[x_8]);
            rqs_00 <= update (update (x_1, x_4, Struct13 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct14
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct13 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct14 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct5) getCRqSlot_00 (Struct4 x_0);
        let x_1 = (rqs_00);
        Struct14 x_2 = (Struct14 {valid : (Bool)'(False), data :
        unpack(0)});
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct14 x_6 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hc)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hc)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hc)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hc)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hd)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hd)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hd)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hd)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'he)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'he)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'he)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'he)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hf)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hf)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hf)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hf)}) : (Struct14 {valid
        : (Bool)'(False), data :
        unpack(0)})))))))))))))))))))))))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(4) x_8 = ((x_6).data);
        Struct5 x_9 = (Struct5 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct13 x_10 = ((x_1)[x_8]);
            rqs_00 <= update (update (x_1, x_4, Struct13 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct14
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct13 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct14 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct7) getWait_00 ();
        let x_1 = (rqs_00);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (((((x_1)[(Bit#(4))'(4'hc)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hc)}) : (((((x_1)[(Bit#(4))'(4'hd)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hd)}) : (((((x_1)[(Bit#(4))'(4'he)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'he)}) : (((((x_1)[(Bit#(4))'(4'hf)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hf)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))))))))))))))))))));
        let x_6 = ?;
        if ((x_2).valid) begin
            Bit#(4) x_3 = ((x_2).data);
            Struct13 x_4 = ((x_1)[x_3]);
            rqs_00 <= update (x_1, x_3, Struct13 {m_status :
            (Bit#(2))'(2'h3), m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul,
            m_msg : (x_4).m_msg, m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb,
            m_dl_rss_from : (x_4).m_dl_rss_from, m_dl_rss_recv :
            (x_4).m_dl_rss_recv, m_dl_rss : (x_4).m_dl_rss});
            Struct4 x_5 = (Struct4 {r_id : x_3, r_msg : (x_4).m_msg,
            r_msg_from : (x_4).m_qidx});
            x_6 = Struct7 {valid : (Bool)'(True), data : x_5};
        end else begin
            x_6 = Struct7 {valid : (Bool)'(False), data : unpack(0)};
        end
        return x_6;
    endmethod

    method Action registerUL_00 (Struct18 x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_00 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_00 (Struct19 x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_00 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(4)) getULImm_00 (Struct1 x_0);
        let x_1 = (rqs_00);
        Struct14 x_2 = (Struct14 {valid : (Bool)'(False), data :
        unpack(0)});
        when ((x_2).valid, noAction);
        Bit#(4) x_3 = ((x_2).data);
        rqs_00 <= update (x_1, x_3, Struct13 {m_status : (Bit#(2))'(2'h3),
        m_next : Struct14 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul
        : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0), m_rsb :
        (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
        m_dl_rss : unpack(0)});
        return x_3;
    endmethod

    method ActionValue#(Bit#(4)) getULCount_00 ();
        let x_1 = (rqs_00);
        Bit#(4) x_2 = ((Bit#(4))'(4'h0));
        return x_2;
    endmethod

    method Action transferUpDown_00 (Struct22 x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_00 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(4)) findUL_00 (Bit#(64) x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = (unpack(0));
        return x_2;
    endmethod

    method ActionValue#(Bit#(4)) findDL_00 (Bit#(64) x_0);
        let x_1 = (rqs_00);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h0)) : (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h1)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h2)) : (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h3)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hb)) : (((((((x_1)[(Bit#(4))'(4'hc)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hc)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hc)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hc)) : (((((((x_1)[(Bit#(4))'(4'hd)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hd)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hd)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hd)) : (((((((x_1)[(Bit#(4))'(4'he)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'he)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'he)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'he)) : (((((((x_1)[(Bit#(4))'(4'hf)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hf)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hf)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hf)) :
        (unpack(0))))))))))))))))))))))))))))))))));
        return x_2;
    endmethod

    method Action releaseMSHR_00 (Bit#(4) x_0);
        let x_1 = (rqs_00);
        Struct13 x_2 = ((x_1)[x_0]);
        Vector#(16, Struct13) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(4) x_4 = (((x_2).m_next).data);
            Struct13 x_5 = ((x_1)[x_4]);
            Vector#(16, Struct13) x_6 = (update (x_3, x_4, Struct13 {m_status
            : (Bit#(2))'(2'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_00 <= x_7;
    endmethod

    method Action addRs_00 (Struct6 x_0);
        let x_1 = (rqs_00);
        Bit#(64) x_2 = (((x_0).r_dl_msg).addr);
        Bit#(4) x_3 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h0)) : (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h1)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h2)) : (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h3)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'hb)) : (((((((x_1)[(Bit#(4))'(4'hc)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hc)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hc)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'hc)) : (((((((x_1)[(Bit#(4))'(4'hd)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hd)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hd)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'hd)) : (((((((x_1)[(Bit#(4))'(4'he)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'he)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'he)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'he)) : (((((((x_1)[(Bit#(4))'(4'hf)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hf)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hf)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'hf)) :
        (unpack(0))))))))))))))))))))))))))))))))));
        Struct13 x_4 = ((x_1)[x_3]);
        Struct13 x_5 = (Struct13 {m_status : (x_4).m_status, m_next :
        (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg, m_qidx :
        (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : ((x_4).m_dl_rss_recv) |
        (((Bit#(2))'(2'h1)) << ((x_0).r_dl_midx)), m_dl_rss : update
        ((x_4).m_dl_rss, (x_0).r_dl_midx, (x_0).r_dl_msg)});
        rqs_00 <= update (x_1, x_3, x_5);
    endmethod

    method ActionValue#(Struct8) getRsReady_00 ();
        let x_1 = (rqs_00);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h0)) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h1)) :
        (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h2)) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h3)) :
        (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h4)) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h5)) :
        (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h6)) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h7)) :
        (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h8)) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h9)) :
        (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'ha)) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'hb)) :
        (((((((x_1)[(Bit#(4))'(4'hc)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'hc)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'hc)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'hc)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'hc)) :
        (((((((x_1)[(Bit#(4))'(4'hd)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'hd)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'hd)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'hd)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'hd)) :
        (((((((x_1)[(Bit#(4))'(4'he)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'he)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'he)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'he)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'he)) :
        (((((((x_1)[(Bit#(4))'(4'hf)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'hf)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'hf)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'hf)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'hf)) :
        (unpack(0))))))))))))))))))))))))))))))))));
        Struct13 x_3 = ((x_1)[x_2]);
        Struct8 x_4 = (Struct8 {r_id : x_2, r_addr :
        ((x_3).m_msg).addr});
        return x_4;
    endmethod
endmodule

interface Module35;
    method Action enq_fifoCRqInput000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput000 ();
endinterface

module mkModule35 (Module35);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifoCRqInput000 (Struct2 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module36;
    method Action enq_fifoCRsInput000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRsInput000 ();
endinterface

module mkModule36 (Module36);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifoCRsInput000 (Struct2 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifoCRsInput000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module37;
    method Action enq_fifoInput000 (Struct3 x_0);
    method ActionValue#(Struct3) deq_fifoInput000 ();
endinterface

module mkModule37 (Module37);
    FIFOF#(Struct3) pff <- mkFIFOF();

    method Action enq_fifoInput000 (Struct3 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct3) deq_fifoInput000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module38;
    method Action enq_fifoI2L000 (Struct3 x_0);
    method ActionValue#(Struct3) deq_fifoI2L000 ();
endinterface

module mkModule38 (Module38);
    FIFOF#(Struct3) pff <- mkFIFOF();

    method Action enq_fifoI2L000 (Struct3 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct3) deq_fifoI2L000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module39;
    method Action enq_fifoL2E000 (Struct42 x_0);
    method ActionValue#(Struct42) deq_fifoL2E000 ();
endinterface

module mkModule39 (Module39);
    FIFOF#(Struct42) pff <- mkFIFOF();

    method Action enq_fifoL2E000 (Struct42 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct42) deq_fifoL2E000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module40;
    method Action enq_fifo0000 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0000 ();
endinterface

module mkModule40 (Module40);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo0000 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo0000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module41;
    method Action enq_fifo0001 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0001 ();
endinterface

module mkModule41 (Module41);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo0001 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo0001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module42;
    method Action enq_fifo0002 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0002 ();
endinterface

module mkModule42 (Module42);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo0002 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo0002 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module43;
    method Action enq_cp_1__000 (Struct44 x_0);
    method ActionValue#(Struct44) deq_cp_1__000 ();
endinterface

module mkModule43 (Module43);
    FIFOF#(Struct44) pff <- mkPipelineFIFOF();

    method Action enq_cp_1__000 (Struct44 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct44) deq_cp_1__000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module44;
    method Action enq_cp_2__000 (Struct45 x_0);
    method ActionValue#(Struct45) deq_cp_2__000 ();
endinterface

module mkModule44 (Module44);
    FIFOF#(Struct45) pff <- mkPipelineFIFOF();

    method Action enq_cp_2__000 (Struct45 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct45) deq_cp_2__000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module45;
    method Action rdReq_infoRam__000__7 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__7 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__7 ();
endinterface

module mkModule45 (Module45);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h7, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__7 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__7 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__7 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module46;
    method Action rdReq_infoRam__000__6 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__6 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__6 ();
endinterface

module mkModule46 (Module46);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h6, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__6 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__6 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__6 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module47;
    method Action rdReq_infoRam__000__5 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__5 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__5 ();
endinterface

module mkModule47 (Module47);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h5, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__5 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__5 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__5 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module48;
    method Action rdReq_infoRam__000__4 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__4 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__4 ();
endinterface

module mkModule48 (Module48);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h4, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__4 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__4 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__4 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module49;
    method Action rdReq_infoRam__000__3 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__3 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__3 ();
endinterface

module mkModule49 (Module49);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h3, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__3 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__3 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module50;
    method Action rdReq_infoRam__000__2 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__2 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__2 ();
endinterface

module mkModule50 (Module50);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h2, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__2 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__2 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module51;
    method Action rdReq_infoRam__000__1 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__1 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__1 ();
endinterface

module mkModule51 (Module51);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h1, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__1 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__1 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module52;
    method Action rdReq_infoRam__000__0 (Bit#(9) x_0);
    method Action wrReq_infoRam__000__0 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__000__0 ();
endinterface

module mkModule52 (Module52);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h0, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__000__0 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__000__0 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__000__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module53;
    method Action rdReq_edirRam__000__3 (Bit#(9) x_0);
    method Action wrReq_edirRam__000__3 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__000__3 ();
endinterface

module mkModule53 (Module53);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h3, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__000__3 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__000__3 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__000__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module54;
    method Action rdReq_edirRam__000__2 (Bit#(9) x_0);
    method Action wrReq_edirRam__000__2 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__000__2 ();
endinterface

module mkModule54 (Module54);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h2, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__000__2 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__000__2 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__000__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module55;
    method Action rdReq_edirRam__000__1 (Bit#(9) x_0);
    method Action wrReq_edirRam__000__1 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__000__1 ();
endinterface

module mkModule55 (Module55);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h1, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__000__1 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__000__1 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__000__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module56;
    method Action rdReq_edirRam__000__0 (Bit#(9) x_0);
    method Action wrReq_edirRam__000__0 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__000__0 ();
endinterface

module mkModule56 (Module56);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h0, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__000__0 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__000__0 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__000__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module57;
    method Action rdReq_dataRam__000 (Bit#(12) x_0);
    method Action wrReq_dataRam__000 (Struct52 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__000 ();
endinterface

module mkModule57 (Module57);
    RWBramCore#(Bit#(12), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(12)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__000 (Bit#(12) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__000 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__000 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module58;
    method Action rdReq_repRam__000 (Bit#(9) x_0);
    method Action wrReq_repRam__000 (Struct54 x_0);
    method ActionValue#(Vector#(8, Bit#(8))) rdResp_repRam__000 ();
endinterface

module mkModule58 (Module58);
    RWBramCore#(Bit#(9), Vector#(8, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__000 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__000 (Struct54 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(8, Bit#(8))) rdResp_repRam__000 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module59;
    method ActionValue#(Struct13) getMSHR_000 (Bit#(4) x_0);
    method ActionValue#(Struct5) getPRqSlot_000 (Struct4 x_0);
    method ActionValue#(Struct5) getCRqSlot_000 (Struct4 x_0);
    method ActionValue#(Struct7) getWait_000 ();
    method Action registerUL_000 (Struct18 x_0);
    method Action registerDL_000 (Struct19 x_0);
    method ActionValue#(Bit#(4)) getULImm_000 (Struct1 x_0);
    method ActionValue#(Bit#(4)) getULCount_000 ();
    method Action transferUpDown_000 (Struct22 x_0);
    method ActionValue#(Bit#(4)) findUL_000 (Bit#(64) x_0);
    method ActionValue#(Bit#(4)) findDL_000 (Bit#(64) x_0);
    method Action releaseMSHR_000 (Bit#(4) x_0);
    method Action addRs_000 (Struct6 x_0);
    method ActionValue#(Struct8) getRsReady_000 ();
endinterface

module mkModule59
    (Module59);
    Reg#(Vector#(12, Struct13)) rqs_000 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct13) getMSHR_000 (Bit#(4) x_0);
        let x_1 = (rqs_000);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct5) getPRqSlot_000 (Struct4 x_0);
        let x_1 = (rqs_000);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct14 x_6 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(4) x_8 = ((x_6).data);
        Struct5 x_9 = (Struct5 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct13 x_10 = ((x_1)[x_8]);
            rqs_000 <= update (update (x_1, x_4, Struct13 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct14
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct13 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct14 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct5) getCRqSlot_000 (Struct4 x_0);
        let x_1 = (rqs_000);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct14 x_6 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(4) x_8 = ((x_6).data);
        Struct5 x_9 = (Struct5 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct13 x_10 = ((x_1)[x_8]);
            rqs_000 <= update (update (x_1, x_4, Struct13 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct14
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct13 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct14 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct7) getWait_000 ();
        let x_1 = (rqs_000);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))))))))))));
        let x_6 = ?;
        if ((x_2).valid) begin
            Bit#(4) x_3 = ((x_2).data);
            Struct13 x_4 = ((x_1)[x_3]);
            rqs_000 <= update (x_1, x_3, Struct13 {m_status :
            (Bit#(2))'(2'h3), m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul,
            m_msg : (x_4).m_msg, m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb,
            m_dl_rss_from : (x_4).m_dl_rss_from, m_dl_rss_recv :
            (x_4).m_dl_rss_recv, m_dl_rss : (x_4).m_dl_rss});
            Struct4 x_5 = (Struct4 {r_id : x_3, r_msg : (x_4).m_msg,
            r_msg_from : (x_4).m_qidx});
            x_6 = Struct7 {valid : (Bool)'(True), data : x_5};
        end else begin
            x_6 = Struct7 {valid : (Bool)'(False), data : unpack(0)};
        end
        return x_6;
    endmethod

    method Action registerUL_000 (Struct18 x_0);
        let x_1 = (rqs_000);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_000 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_000 (Struct19 x_0);
        let x_1 = (rqs_000);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_000 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(4)) getULImm_000 (Struct1 x_0);
        let x_1 = (rqs_000);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hc)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hd)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'he)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hf)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))));
        when ((x_2).valid, noAction);
        Bit#(4) x_3 = ((x_2).data);
        rqs_000 <= update (x_1, x_3, Struct13 {m_status : (Bit#(2))'(2'h3),
        m_next : Struct14 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul
        : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0), m_rsb :
        (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
        m_dl_rss : unpack(0)});
        return x_3;
    endmethod

    method ActionValue#(Bit#(4)) getULCount_000 ();
        let x_1 = (rqs_000);
        Bit#(4) x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'h5)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + (((((x_1)[(Bit#(4))'(4'h6)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'h7)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + (((((x_1)[(Bit#(4))'(4'h8)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'h9)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + (((((x_1)[(Bit#(4))'(4'ha)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'hb)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + ((Bit#(4))'(4'h0))))))))));
        return x_2;
    endmethod

    method Action transferUpDown_000 (Struct22 x_0);
        let x_1 = (rqs_000);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_000 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(4)) findUL_000 (Bit#(64) x_0);
        let x_1 = (rqs_000);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hb)) : (unpack(0))))))))))))))))));
        return x_2;
    endmethod

    method ActionValue#(Bit#(4)) findDL_000 (Bit#(64) x_0);
        let x_1 = (rqs_000);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h0)) : (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h1)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h2)) : (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h3)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hb)) : (unpack(0))))))))))))))))))))))))));
        return x_2;
    endmethod

    method Action releaseMSHR_000 (Bit#(4) x_0);
        let x_1 = (rqs_000);
        Struct13 x_2 = ((x_1)[x_0]);
        Vector#(12, Struct13) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(4) x_4 = (((x_2).m_next).data);
            Struct13 x_5 = ((x_1)[x_4]);
            Vector#(12, Struct13) x_6 = (update (x_3, x_4, Struct13 {m_status
            : (Bit#(2))'(2'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_000 <= x_7;
    endmethod

    method Action addRs_000 (Struct6 x_0);
        let x_1 = (rqs_000);
        Bit#(64) x_2 = (((x_0).r_dl_msg).addr);
        Bit#(4) x_3 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h0)) : (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h1)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h2)) : (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h3)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'hb)) : (unpack(0))))))))))))))))))))))))));
        Struct13 x_4 = ((x_1)[x_3]);
        Struct13 x_5 = (Struct13 {m_status : (x_4).m_status, m_next :
        (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg, m_qidx :
        (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : ((x_4).m_dl_rss_recv) |
        (((Bit#(2))'(2'h1)) << ((x_0).r_dl_midx)), m_dl_rss : update
        ((x_4).m_dl_rss, (x_0).r_dl_midx, (x_0).r_dl_msg)});
        rqs_000 <= update (x_1, x_3, x_5);
    endmethod

    method ActionValue#(Struct8) getRsReady_000 ();
        let x_1 = (rqs_000);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h0)) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h1)) :
        (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h2)) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h3)) :
        (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h4)) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h5)) :
        (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h6)) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h7)) :
        (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h8)) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h9)) :
        (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'ha)) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'hb)) :
        (unpack(0))))))))))))))))))))))))));
        Struct13 x_3 = ((x_1)[x_2]);
        Struct8 x_4 = (Struct8 {r_id : x_2, r_addr :
        ((x_3).m_msg).addr});
        return x_4;
    endmethod
endmodule

interface Module60;
    method Action enq_fifoInput0000 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoInput0000 ();
endinterface

module mkModule60 (Module60);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoInput0000 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoInput0000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module61;
    method Action enq_fifoI2L0000 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoI2L0000 ();
endinterface

module mkModule61 (Module61);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoI2L0000 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoI2L0000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module62;
    method Action enq_fifoL2E0000 (Struct62 x_0);
    method ActionValue#(Struct62) deq_fifoL2E0000 ();
endinterface

module mkModule62 (Module62);
    FIFOF#(Struct62) pff <- mkFIFOF();

    method Action enq_fifoL2E0000 (Struct62 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct62) deq_fifoL2E0000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module63;
    method Action enq_fifo00000 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00000 ();
endinterface

module mkModule63 (Module63);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00000 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module64;
    method Action enq_fifo00001 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00001 ();
endinterface

module mkModule64 (Module64);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00001 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module65;
    method Action enq_fifo00002 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00002 ();
endinterface

module mkModule65 (Module65);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00002 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00002 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module66;
    method Action enq_fifo000000 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo000000 ();
endinterface

module mkModule66 (Module66);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo000000 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo000000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module67;
    method Action enq_fifo000002 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo000002 ();
endinterface

module mkModule67 (Module67);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo000002 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo000002 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module68;
    method Action enq_cp_1__0000 (Struct68 x_0);
    method ActionValue#(Struct68) deq_cp_1__0000 ();
endinterface

module mkModule68 (Module68);
    FIFOF#(Struct68) pff <- mkPipelineFIFOF();

    method Action enq_cp_1__0000 (Struct68 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct68) deq_cp_1__0000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module69;
    method Action enq_cp_2__0000 (Struct69 x_0);
    method ActionValue#(Struct69) deq_cp_2__0000 ();
endinterface

module mkModule69 (Module69);
    FIFOF#(Struct69) pff <- mkPipelineFIFOF();

    method Action enq_cp_2__0000 (Struct69 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct69) deq_cp_2__0000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module70;
    method Action rdReq_infoRam__0000__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__0000__3 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0000__3 ();
endinterface

module mkModule70 (Module70);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h3, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0000__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0000__3 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0000__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module71;
    method Action rdReq_infoRam__0000__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__0000__2 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0000__2 ();
endinterface

module mkModule71 (Module71);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h2, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0000__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0000__2 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0000__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module72;
    method Action rdReq_infoRam__0000__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__0000__1 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0000__1 ();
endinterface

module mkModule72 (Module72);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h1, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0000__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0000__1 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0000__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module73;
    method Action rdReq_infoRam__0000__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__0000__0 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0000__0 ();
endinterface

module mkModule73 (Module73);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h0, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0000__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0000__0 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0000__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module74;
    method Action rdReq_dataRam__0000 (Bit#(10) x_0);
    method Action wrReq_dataRam__0000 (Struct73 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0000 ();
endinterface

module mkModule74 (Module74);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__0000 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__0000 (Struct73 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0000 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module75;
    method Action rdReq_repRam__0000 (Bit#(8) x_0);
    method Action wrReq_repRam__0000 (Struct76 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0000 ();
endinterface

module mkModule75 (Module75);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h0, 8'h0, 8'h0, 8'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__0000 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__0000 (Struct76 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0000 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module76;
    method ActionValue#(Struct63) getMSHR_0000 (Bit#(3) x_0);
    method ActionValue#(Struct57) getPRqSlot_0000 (Struct56 x_0);
    method ActionValue#(Struct57) getCRqSlot_0000 (Struct56 x_0);
    method ActionValue#(Struct58) getWait_0000 ();
    method Action registerUL_0000 (Struct65 x_0);
    method Action registerDL_0000 (Struct77 x_0);
    method ActionValue#(Bit#(3)) getULImm_0000 (Struct1 x_0);
    method ActionValue#(Bit#(3)) getULCount_0000 ();
    method Action transferUpDown_0000 (Struct78 x_0);
    method ActionValue#(Bit#(3)) findUL_0000 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) findDL_0000 (Bit#(64) x_0);
    method Action releaseMSHR_0000 (Bit#(3) x_0);
    method Action addRs_0000 (Struct6 x_0);
    method ActionValue#(Struct59) getRsReady_0000 ();
endinterface

module mkModule76
    (Module76);
    Reg#(Vector#(6, Struct63)) rqs_0000 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct63) getMSHR_0000 (Bit#(3) x_0);
        let x_1 = (rqs_0000);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct57) getPRqSlot_0000 (Struct56 x_0);
        let x_1 = (rqs_0000);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0000 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct57) getCRqSlot_0000 (Struct56 x_0);
        let x_1 = (rqs_0000);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0000 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct58) getWait_0000 ();
        let x_1 = (rqs_0000);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        let x_6 = ?;
        if ((x_2).valid) begin
            Bit#(3) x_3 = ((x_2).data);
            Struct63 x_4 = ((x_1)[x_3]);
            rqs_0000 <= update (x_1, x_3, Struct63 {m_status :
            (Bit#(2))'(2'h3), m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul,
            m_msg : (x_4).m_msg, m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb,
            m_dl_rss_from : (x_4).m_dl_rss_from, m_dl_rss_recv :
            (x_4).m_dl_rss_recv, m_dl_rss : (x_4).m_dl_rss});
            Struct56 x_5 = (Struct56 {r_id : x_3, r_msg : (x_4).m_msg,
            r_msg_from : (x_4).m_qidx});
            x_6 = Struct58 {valid : (Bool)'(True), data : x_5};
        end else begin
            x_6 = Struct58 {valid : (Bool)'(False), data : unpack(0)};
        end
        return x_6;
    endmethod

    method Action registerUL_0000 (Struct65 x_0);
        let x_1 = (rqs_0000);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_0000 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_0000 (Struct77 x_0);
        let x_1 = (rqs_0000);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0000 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) getULImm_0000 (Struct1 x_0);
        let x_1 = (rqs_0000);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h6)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h7)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        rqs_0000 <= update (x_1, x_3, Struct63 {m_status : (Bit#(2))'(2'h3),
        m_next : Struct10 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul
        : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0), m_rsb :
        (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
        m_dl_rss : unpack(0)});
        return x_3;
    endmethod

    method ActionValue#(Bit#(3)) getULCount_0000 ();
        let x_1 = (rqs_0000);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h3)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + (((((x_1)[(Bit#(3))'(3'h4)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h5)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + ((Bit#(3))'(3'h0))))));
        return x_2;
    endmethod

    method Action transferUpDown_0000 (Struct78 x_0);
        let x_1 = (rqs_0000);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0000 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) findUL_0000 (Bit#(64) x_0);
        let x_1 = (rqs_0000);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))));
        return x_2;
    endmethod

    method ActionValue#(Bit#(3)) findDL_0000 (Bit#(64) x_0);
        let x_1 = (rqs_0000);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        return x_2;
    endmethod

    method Action releaseMSHR_0000 (Bit#(3) x_0);
        let x_1 = (rqs_0000);
        Struct63 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct63) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct63 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct63) x_6 = (update (x_3, x_4, Struct63 {m_status
            : (Bit#(2))'(2'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_0000 <= x_7;
    endmethod

    method Action addRs_0000 (Struct6 x_0);
        let x_1 = (rqs_0000);
        Bit#(64) x_2 = (((x_0).r_dl_msg).addr);
        Bit#(3) x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        Struct63 x_4 = ((x_1)[x_3]);
        Struct63 x_5 = (Struct63 {m_status : (x_4).m_status, m_next :
        (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg, m_qidx :
        (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : ((x_4).m_dl_rss_recv) |
        (((Bit#(2))'(2'h1)) << ((x_0).r_dl_midx)), m_dl_rss : update
        ((x_4).m_dl_rss, (x_0).r_dl_midx, (x_0).r_dl_msg)});
        rqs_0000 <= update (x_1, x_3, x_5);
    endmethod

    method ActionValue#(Struct59) getRsReady_0000 ();
        let x_1 = (rqs_0000);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h0)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h1)) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h2)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h3)) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h4)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h5)) :
        (unpack(0))))))))))))));
        Struct63 x_3 = ((x_1)[x_2]);
        Struct59 x_4 = (Struct59 {r_id : x_2, r_addr :
        ((x_3).m_msg).addr});
        return x_4;
    endmethod
endmodule

interface Module77;
    method Action enq_fifoInput0001 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoInput0001 ();
endinterface

module mkModule77 (Module77);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoInput0001 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoInput0001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module78;
    method Action enq_fifoI2L0001 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoI2L0001 ();
endinterface

module mkModule78 (Module78);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoI2L0001 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoI2L0001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module79;
    method Action enq_fifoL2E0001 (Struct62 x_0);
    method ActionValue#(Struct62) deq_fifoL2E0001 ();
endinterface

module mkModule79 (Module79);
    FIFOF#(Struct62) pff <- mkFIFOF();

    method Action enq_fifoL2E0001 (Struct62 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct62) deq_fifoL2E0001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module80;
    method Action enq_fifo00010 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00010 ();
endinterface

module mkModule80 (Module80);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00010 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00010 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module81;
    method Action enq_fifo00011 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00011 ();
endinterface

module mkModule81 (Module81);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00011 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00011 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module82;
    method Action enq_fifo00012 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00012 ();
endinterface

module mkModule82 (Module82);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00012 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00012 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module83;
    method Action enq_fifo000100 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo000100 ();
endinterface

module mkModule83 (Module83);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo000100 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo000100 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module84;
    method Action enq_fifo000102 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo000102 ();
endinterface

module mkModule84 (Module84);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo000102 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo000102 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module85;
    method Action enq_cp_1__0001 (Struct68 x_0);
    method ActionValue#(Struct68) deq_cp_1__0001 ();
endinterface

module mkModule85 (Module85);
    FIFOF#(Struct68) pff <- mkPipelineFIFOF();

    method Action enq_cp_1__0001 (Struct68 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct68) deq_cp_1__0001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module86;
    method Action enq_cp_2__0001 (Struct69 x_0);
    method ActionValue#(Struct69) deq_cp_2__0001 ();
endinterface

module mkModule86 (Module86);
    FIFOF#(Struct69) pff <- mkPipelineFIFOF();

    method Action enq_cp_2__0001 (Struct69 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct69) deq_cp_2__0001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module87;
    method Action rdReq_infoRam__0001__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__0001__3 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0001__3 ();
endinterface

module mkModule87 (Module87);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h3, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0001__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0001__3 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0001__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module88;
    method Action rdReq_infoRam__0001__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__0001__2 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0001__2 ();
endinterface

module mkModule88 (Module88);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h2, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0001__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0001__2 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0001__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module89;
    method Action rdReq_infoRam__0001__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__0001__1 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0001__1 ();
endinterface

module mkModule89 (Module89);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h1, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0001__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0001__1 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0001__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module90;
    method Action rdReq_infoRam__0001__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__0001__0 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0001__0 ();
endinterface

module mkModule90 (Module90);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h0, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0001__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0001__0 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0001__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module91;
    method Action rdReq_dataRam__0001 (Bit#(10) x_0);
    method Action wrReq_dataRam__0001 (Struct73 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0001 ();
endinterface

module mkModule91 (Module91);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__0001 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__0001 (Struct73 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0001 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module92;
    method Action rdReq_repRam__0001 (Bit#(8) x_0);
    method Action wrReq_repRam__0001 (Struct76 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0001 ();
endinterface

module mkModule92 (Module92);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h0, 8'h0, 8'h0, 8'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__0001 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__0001 (Struct76 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0001 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module93;
    method ActionValue#(Struct63) getMSHR_0001 (Bit#(3) x_0);
    method ActionValue#(Struct57) getPRqSlot_0001 (Struct56 x_0);
    method ActionValue#(Struct57) getCRqSlot_0001 (Struct56 x_0);
    method ActionValue#(Struct58) getWait_0001 ();
    method Action registerUL_0001 (Struct65 x_0);
    method Action registerDL_0001 (Struct77 x_0);
    method ActionValue#(Bit#(3)) getULImm_0001 (Struct1 x_0);
    method ActionValue#(Bit#(3)) getULCount_0001 ();
    method Action transferUpDown_0001 (Struct78 x_0);
    method ActionValue#(Bit#(3)) findUL_0001 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) findDL_0001 (Bit#(64) x_0);
    method Action releaseMSHR_0001 (Bit#(3) x_0);
    method Action addRs_0001 (Struct6 x_0);
    method ActionValue#(Struct59) getRsReady_0001 ();
endinterface

module mkModule93
    (Module93);
    Reg#(Vector#(6, Struct63)) rqs_0001 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct63) getMSHR_0001 (Bit#(3) x_0);
        let x_1 = (rqs_0001);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct57) getPRqSlot_0001 (Struct56 x_0);
        let x_1 = (rqs_0001);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0001 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct57) getCRqSlot_0001 (Struct56 x_0);
        let x_1 = (rqs_0001);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0001 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct58) getWait_0001 ();
        let x_1 = (rqs_0001);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        let x_6 = ?;
        if ((x_2).valid) begin
            Bit#(3) x_3 = ((x_2).data);
            Struct63 x_4 = ((x_1)[x_3]);
            rqs_0001 <= update (x_1, x_3, Struct63 {m_status :
            (Bit#(2))'(2'h3), m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul,
            m_msg : (x_4).m_msg, m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb,
            m_dl_rss_from : (x_4).m_dl_rss_from, m_dl_rss_recv :
            (x_4).m_dl_rss_recv, m_dl_rss : (x_4).m_dl_rss});
            Struct56 x_5 = (Struct56 {r_id : x_3, r_msg : (x_4).m_msg,
            r_msg_from : (x_4).m_qidx});
            x_6 = Struct58 {valid : (Bool)'(True), data : x_5};
        end else begin
            x_6 = Struct58 {valid : (Bool)'(False), data : unpack(0)};
        end
        return x_6;
    endmethod

    method Action registerUL_0001 (Struct65 x_0);
        let x_1 = (rqs_0001);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_0001 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_0001 (Struct77 x_0);
        let x_1 = (rqs_0001);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0001 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) getULImm_0001 (Struct1 x_0);
        let x_1 = (rqs_0001);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h6)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h7)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        rqs_0001 <= update (x_1, x_3, Struct63 {m_status : (Bit#(2))'(2'h3),
        m_next : Struct10 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul
        : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0), m_rsb :
        (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
        m_dl_rss : unpack(0)});
        return x_3;
    endmethod

    method ActionValue#(Bit#(3)) getULCount_0001 ();
        let x_1 = (rqs_0001);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h3)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + (((((x_1)[(Bit#(3))'(3'h4)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h5)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + ((Bit#(3))'(3'h0))))));
        return x_2;
    endmethod

    method Action transferUpDown_0001 (Struct78 x_0);
        let x_1 = (rqs_0001);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0001 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) findUL_0001 (Bit#(64) x_0);
        let x_1 = (rqs_0001);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))));
        return x_2;
    endmethod

    method ActionValue#(Bit#(3)) findDL_0001 (Bit#(64) x_0);
        let x_1 = (rqs_0001);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        return x_2;
    endmethod

    method Action releaseMSHR_0001 (Bit#(3) x_0);
        let x_1 = (rqs_0001);
        Struct63 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct63) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct63 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct63) x_6 = (update (x_3, x_4, Struct63 {m_status
            : (Bit#(2))'(2'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_0001 <= x_7;
    endmethod

    method Action addRs_0001 (Struct6 x_0);
        let x_1 = (rqs_0001);
        Bit#(64) x_2 = (((x_0).r_dl_msg).addr);
        Bit#(3) x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        Struct63 x_4 = ((x_1)[x_3]);
        Struct63 x_5 = (Struct63 {m_status : (x_4).m_status, m_next :
        (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg, m_qidx :
        (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : ((x_4).m_dl_rss_recv) |
        (((Bit#(2))'(2'h1)) << ((x_0).r_dl_midx)), m_dl_rss : update
        ((x_4).m_dl_rss, (x_0).r_dl_midx, (x_0).r_dl_msg)});
        rqs_0001 <= update (x_1, x_3, x_5);
    endmethod

    method ActionValue#(Struct59) getRsReady_0001 ();
        let x_1 = (rqs_0001);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h0)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h1)) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h2)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h3)) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h4)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h5)) :
        (unpack(0))))))))))))));
        Struct63 x_3 = ((x_1)[x_2]);
        Struct59 x_4 = (Struct59 {r_id : x_2, r_addr :
        ((x_3).m_msg).addr});
        return x_4;
    endmethod
endmodule

interface Module94;
    method Action enq_fifoCRqInput001 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRqInput001 ();
endinterface

module mkModule94 (Module94);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifoCRqInput001 (Struct2 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifoCRqInput001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module95;
    method Action enq_fifoCRsInput001 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifoCRsInput001 ();
endinterface

module mkModule95 (Module95);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifoCRsInput001 (Struct2 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifoCRsInput001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module96;
    method Action enq_fifoInput001 (Struct3 x_0);
    method ActionValue#(Struct3) deq_fifoInput001 ();
endinterface

module mkModule96 (Module96);
    FIFOF#(Struct3) pff <- mkFIFOF();

    method Action enq_fifoInput001 (Struct3 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct3) deq_fifoInput001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module97;
    method Action enq_fifoI2L001 (Struct3 x_0);
    method ActionValue#(Struct3) deq_fifoI2L001 ();
endinterface

module mkModule97 (Module97);
    FIFOF#(Struct3) pff <- mkFIFOF();

    method Action enq_fifoI2L001 (Struct3 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct3) deq_fifoI2L001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module98;
    method Action enq_fifoL2E001 (Struct42 x_0);
    method ActionValue#(Struct42) deq_fifoL2E001 ();
endinterface

module mkModule98 (Module98);
    FIFOF#(Struct42) pff <- mkFIFOF();

    method Action enq_fifoL2E001 (Struct42 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct42) deq_fifoL2E001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module99;
    method Action enq_fifo0010 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0010 ();
endinterface

module mkModule99 (Module99);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo0010 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo0010 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module100;
    method Action enq_fifo0011 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0011 ();
endinterface

module mkModule100 (Module100);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo0011 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo0011 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module101;
    method Action enq_fifo0012 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo0012 ();
endinterface

module mkModule101 (Module101);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo0012 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo0012 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module102;
    method Action enq_cp_1__001 (Struct44 x_0);
    method ActionValue#(Struct44) deq_cp_1__001 ();
endinterface

module mkModule102 (Module102);
    FIFOF#(Struct44) pff <- mkPipelineFIFOF();

    method Action enq_cp_1__001 (Struct44 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct44) deq_cp_1__001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module103;
    method Action enq_cp_2__001 (Struct45 x_0);
    method ActionValue#(Struct45) deq_cp_2__001 ();
endinterface

module mkModule103 (Module103);
    FIFOF#(Struct45) pff <- mkPipelineFIFOF();

    method Action enq_cp_2__001 (Struct45 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct45) deq_cp_2__001 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module104;
    method Action rdReq_infoRam__001__7 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__7 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__7 ();
endinterface

module mkModule104 (Module104);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h7, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__7 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__7 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__7 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module105;
    method Action rdReq_infoRam__001__6 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__6 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__6 ();
endinterface

module mkModule105 (Module105);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h6, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__6 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__6 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__6 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module106;
    method Action rdReq_infoRam__001__5 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__5 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__5 ();
endinterface

module mkModule106 (Module106);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h5, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__5 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__5 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__5 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module107;
    method Action rdReq_infoRam__001__4 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__4 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__4 ();
endinterface

module mkModule107 (Module107);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h4, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__4 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__4 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__4 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module108;
    method Action rdReq_infoRam__001__3 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__3 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__3 ();
endinterface

module mkModule108 (Module108);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h3, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__3 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__3 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module109;
    method Action rdReq_infoRam__001__2 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__2 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__2 ();
endinterface

module mkModule109 (Module109);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h2, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__2 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__2 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module110;
    method Action rdReq_infoRam__001__1 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__1 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__1 ();
endinterface

module mkModule110 (Module110);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h1, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__1 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__1 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module111;
    method Action rdReq_infoRam__001__0 (Bit#(9) x_0);
    method Action wrReq_infoRam__001__0 (Struct50 x_0);
    method ActionValue#(Struct46) rdResp_infoRam__001__0 ();
endinterface

module mkModule111 (Module111);
    RWBramCore#(Bit#(9), Struct46) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct46 {tag: 50'h0, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__001__0 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__001__0 (Struct50 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct46) rdResp_infoRam__001__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module112;
    method Action rdReq_edirRam__001__3 (Bit#(9) x_0);
    method Action wrReq_edirRam__001__3 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__001__3 ();
endinterface

module mkModule112 (Module112);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h3, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__001__3 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__001__3 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__001__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module113;
    method Action rdReq_edirRam__001__2 (Bit#(9) x_0);
    method Action wrReq_edirRam__001__2 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__001__2 ();
endinterface

module mkModule113 (Module113);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h2, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__001__2 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__001__2 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__001__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module114;
    method Action rdReq_edirRam__001__1 (Bit#(9) x_0);
    method Action wrReq_edirRam__001__1 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__001__1 ();
endinterface

module mkModule114 (Module114);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h1, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__001__1 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__001__1 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__001__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module115;
    method Action rdReq_edirRam__001__0 (Bit#(9) x_0);
    method Action wrReq_edirRam__001__0 (Struct53 x_0);
    method ActionValue#(Struct48) rdResp_edirRam__001__0 ();
endinterface

module mkModule115 (Module115);
    RWBramCore#(Bit#(9), Struct48) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct48 {tag: 50'h0, value: Struct32 {mesi_edir_st: 3'h1, mesi_edir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_edirRam__001__0 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_edirRam__001__0 (Struct53 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct48) rdResp_edirRam__001__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module116;
    method Action rdReq_dataRam__001 (Bit#(12) x_0);
    method Action wrReq_dataRam__001 (Struct52 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__001 ();
endinterface

module mkModule116 (Module116);
    RWBramCore#(Bit#(12), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(12)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__001 (Bit#(12) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__001 (Struct52 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__001 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module117;
    method Action rdReq_repRam__001 (Bit#(9) x_0);
    method Action wrReq_repRam__001 (Struct54 x_0);
    method ActionValue#(Vector#(8, Bit#(8))) rdResp_repRam__001 ();
endinterface

module mkModule117 (Module117);
    RWBramCore#(Bit#(9), Vector#(8, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(9)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0, 8'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__001 (Bit#(9) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__001 (Struct54 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(8, Bit#(8))) rdResp_repRam__001 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module118;
    method ActionValue#(Struct13) getMSHR_001 (Bit#(4) x_0);
    method ActionValue#(Struct5) getPRqSlot_001 (Struct4 x_0);
    method ActionValue#(Struct5) getCRqSlot_001 (Struct4 x_0);
    method ActionValue#(Struct7) getWait_001 ();
    method Action registerUL_001 (Struct18 x_0);
    method Action registerDL_001 (Struct19 x_0);
    method ActionValue#(Bit#(4)) getULImm_001 (Struct1 x_0);
    method ActionValue#(Bit#(4)) getULCount_001 ();
    method Action transferUpDown_001 (Struct22 x_0);
    method ActionValue#(Bit#(4)) findUL_001 (Bit#(64) x_0);
    method ActionValue#(Bit#(4)) findDL_001 (Bit#(64) x_0);
    method Action releaseMSHR_001 (Bit#(4) x_0);
    method Action addRs_001 (Struct6 x_0);
    method ActionValue#(Struct8) getRsReady_001 ();
endinterface

module mkModule118
    (Module118);
    Reg#(Vector#(12, Struct13)) rqs_001 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct13) getMSHR_001 (Bit#(4) x_0);
        let x_1 = (rqs_001);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct5) getPRqSlot_001 (Struct4 x_0);
        let x_1 = (rqs_001);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct14 x_6 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(4) x_8 = ((x_6).data);
        Struct5 x_9 = (Struct5 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct13 x_10 = ((x_1)[x_8]);
            rqs_001 <= update (update (x_1, x_4, Struct13 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct14
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct13 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct14 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct5) getCRqSlot_001 (Struct4 x_0);
        let x_1 = (rqs_001);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(4) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct14 x_6 = ((((! ((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h0)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h1)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h2)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h3)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h4)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h5)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h6)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h6)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h7)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h7)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h8)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h8)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'h9)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'h9)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'ha)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'ha)}) : ((((!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(4))'(4'hb)]).m_next).valid))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_5)) ? (Struct14
        {valid : (Bool)'(True), data : (Bit#(4))'(4'hb)}) : (Struct14 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))))))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(4) x_8 = ((x_6).data);
        Struct5 x_9 = (Struct5 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct13 x_10 = ((x_1)[x_8]);
            rqs_001 <= update (update (x_1, x_4, Struct13 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct14
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct13 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct14 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct7) getWait_001 ();
        let x_1 = (rqs_001);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h0)}) : (((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h1)}) : (((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h2)}) : (((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h3)}) : (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h4)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h5)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h6)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h7)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))))))))))));
        let x_6 = ?;
        if ((x_2).valid) begin
            Bit#(4) x_3 = ((x_2).data);
            Struct13 x_4 = ((x_1)[x_3]);
            rqs_001 <= update (x_1, x_3, Struct13 {m_status :
            (Bit#(2))'(2'h3), m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul,
            m_msg : (x_4).m_msg, m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb,
            m_dl_rss_from : (x_4).m_dl_rss_from, m_dl_rss_recv :
            (x_4).m_dl_rss_recv, m_dl_rss : (x_4).m_dl_rss});
            Struct4 x_5 = (Struct4 {r_id : x_3, r_msg : (x_4).m_msg,
            r_msg_from : (x_4).m_qidx});
            x_6 = Struct7 {valid : (Bool)'(True), data : x_5};
        end else begin
            x_6 = Struct7 {valid : (Bool)'(False), data : unpack(0)};
        end
        return x_6;
    endmethod

    method Action registerUL_001 (Struct18 x_0);
        let x_1 = (rqs_001);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_001 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_001 (Struct19 x_0);
        let x_1 = (rqs_001);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_001 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(4)) getULImm_001 (Struct1 x_0);
        let x_1 = (rqs_001);
        Struct14 x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h8)}) : (((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'h9)}) : (((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'ha)}) : (((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hb)}) : (((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hc)}) : (((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hd)}) : (((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'he)}) : (((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct14 {valid : (Bool)'(True), data :
        (Bit#(4))'(4'hf)}) : (Struct14 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))))))));
        when ((x_2).valid, noAction);
        Bit#(4) x_3 = ((x_2).data);
        rqs_001 <= update (x_1, x_3, Struct13 {m_status : (Bit#(2))'(2'h3),
        m_next : Struct14 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul
        : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0), m_rsb :
        (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
        m_dl_rss : unpack(0)});
        return x_3;
    endmethod

    method ActionValue#(Bit#(4)) getULCount_001 ();
        let x_1 = (rqs_001);
        Bit#(4) x_2 = (((((x_1)[(Bit#(4))'(4'h4)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'h5)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + (((((x_1)[(Bit#(4))'(4'h6)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'h7)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + (((((x_1)[(Bit#(4))'(4'h8)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'h9)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + (((((x_1)[(Bit#(4))'(4'ha)]).m_is_ul ?
        ((Bit#(4))'(4'h1)) : ((Bit#(4))'(4'h0)))) +
        (((((x_1)[(Bit#(4))'(4'hb)]).m_is_ul ? ((Bit#(4))'(4'h1)) :
        ((Bit#(4))'(4'h0)))) + ((Bit#(4))'(4'h0))))))))));
        return x_2;
    endmethod

    method Action transferUpDown_001 (Struct22 x_0);
        let x_1 = (rqs_001);
        Bit#(4) x_2 = ((x_0).r_id);
        Struct13 x_3 = ((x_1)[x_2]);
        Struct13 x_4 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_001 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(4)) findUL_001 (Bit#(64) x_0);
        let x_1 = (rqs_001);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul)) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hb)) : (unpack(0))))))))))))))))));
        return x_2;
    endmethod

    method ActionValue#(Bit#(4)) findDL_001 (Bit#(64) x_0);
        let x_1 = (rqs_001);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h0)) : (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h1)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h2)) : (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h3)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_0)) ?
        ((Bit#(4))'(4'hb)) : (unpack(0))))))))))))))))))))))))));
        return x_2;
    endmethod

    method Action releaseMSHR_001 (Bit#(4) x_0);
        let x_1 = (rqs_001);
        Struct13 x_2 = ((x_1)[x_0]);
        Vector#(12, Struct13) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(4) x_4 = (((x_2).m_next).data);
            Struct13 x_5 = ((x_1)[x_4]);
            Vector#(12, Struct13) x_6 = (update (x_3, x_4, Struct13 {m_status
            : (Bit#(2))'(2'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_001 <= x_7;
    endmethod

    method Action addRs_001 (Struct6 x_0);
        let x_1 = (rqs_001);
        Bit#(64) x_2 = (((x_0).r_dl_msg).addr);
        Bit#(4) x_3 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h0)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h0)) : (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h1)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h1)) : (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h2)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h2)) : (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h3)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h3)) : (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h4)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h4)) : (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h5)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h5)) : (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h6)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h6)) : (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h7)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h7)) : (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h8)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h8)) : (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'h9)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'h9)) : (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'ha)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'ha)) : (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        (((((x_1)[(Bit#(4))'(4'hb)]).m_msg).addr) == (x_2)) ?
        ((Bit#(4))'(4'hb)) : (unpack(0))))))))))))))))))))))))));
        Struct13 x_4 = ((x_1)[x_3]);
        Struct13 x_5 = (Struct13 {m_status : (x_4).m_status, m_next :
        (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg, m_qidx :
        (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : ((x_4).m_dl_rss_recv) |
        (((Bit#(2))'(2'h1)) << ((x_0).r_dl_midx)), m_dl_rss : update
        ((x_4).m_dl_rss, (x_0).r_dl_midx, (x_0).r_dl_msg)});
        rqs_001 <= update (x_1, x_3, x_5);
    endmethod

    method ActionValue#(Struct8) getRsReady_001 ();
        let x_1 = (rqs_001);
        Bit#(4) x_2 = (((((((x_1)[(Bit#(4))'(4'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(4))'(4'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h0)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h0)) :
        (((((((x_1)[(Bit#(4))'(4'h1)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h1)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h1)) :
        (((((((x_1)[(Bit#(4))'(4'h2)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h2)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h2)) :
        (((((((x_1)[(Bit#(4))'(4'h3)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h3)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h3)) :
        (((((((x_1)[(Bit#(4))'(4'h4)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h4)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h4)) :
        (((((((x_1)[(Bit#(4))'(4'h5)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h5)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h5)) :
        (((((((x_1)[(Bit#(4))'(4'h6)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h6)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h6)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h6)) :
        (((((((x_1)[(Bit#(4))'(4'h7)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h7)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h7)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h7)) :
        (((((((x_1)[(Bit#(4))'(4'h8)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h8)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h8)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h8)) :
        (((((((x_1)[(Bit#(4))'(4'h9)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'h9)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'h9)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'h9)) :
        (((((((x_1)[(Bit#(4))'(4'ha)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'ha)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'ha)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'ha)) :
        (((((((x_1)[(Bit#(4))'(4'hb)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(4))'(4'hb)]).m_is_ul))) &&
        ((((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(4))'(4'hb)]).m_dl_rss_recv)) ? ((Bit#(4))'(4'hb)) :
        (unpack(0))))))))))))))))))))))))));
        Struct13 x_3 = ((x_1)[x_2]);
        Struct8 x_4 = (Struct8 {r_id : x_2, r_addr :
        ((x_3).m_msg).addr});
        return x_4;
    endmethod
endmodule

interface Module119;
    method Action enq_fifoInput0010 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoInput0010 ();
endinterface

module mkModule119 (Module119);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoInput0010 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoInput0010 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module120;
    method Action enq_fifoI2L0010 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoI2L0010 ();
endinterface

module mkModule120 (Module120);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoI2L0010 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoI2L0010 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module121;
    method Action enq_fifoL2E0010 (Struct62 x_0);
    method ActionValue#(Struct62) deq_fifoL2E0010 ();
endinterface

module mkModule121 (Module121);
    FIFOF#(Struct62) pff <- mkFIFOF();

    method Action enq_fifoL2E0010 (Struct62 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct62) deq_fifoL2E0010 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module122;
    method Action enq_fifo00100 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00100 ();
endinterface

module mkModule122 (Module122);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00100 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00100 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module123;
    method Action enq_fifo00101 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00101 ();
endinterface

module mkModule123 (Module123);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00101 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00101 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module124;
    method Action enq_fifo00102 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00102 ();
endinterface

module mkModule124 (Module124);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00102 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00102 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module125;
    method Action enq_fifo001000 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo001000 ();
endinterface

module mkModule125 (Module125);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo001000 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo001000 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module126;
    method Action enq_fifo001002 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo001002 ();
endinterface

module mkModule126 (Module126);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo001002 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo001002 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module127;
    method Action enq_cp_1__0010 (Struct68 x_0);
    method ActionValue#(Struct68) deq_cp_1__0010 ();
endinterface

module mkModule127 (Module127);
    FIFOF#(Struct68) pff <- mkPipelineFIFOF();

    method Action enq_cp_1__0010 (Struct68 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct68) deq_cp_1__0010 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module128;
    method Action enq_cp_2__0010 (Struct69 x_0);
    method ActionValue#(Struct69) deq_cp_2__0010 ();
endinterface

module mkModule128 (Module128);
    FIFOF#(Struct69) pff <- mkPipelineFIFOF();

    method Action enq_cp_2__0010 (Struct69 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct69) deq_cp_2__0010 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module129;
    method Action rdReq_infoRam__0010__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__0010__3 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0010__3 ();
endinterface

module mkModule129 (Module129);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h3, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0010__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0010__3 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0010__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module130;
    method Action rdReq_infoRam__0010__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__0010__2 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0010__2 ();
endinterface

module mkModule130 (Module130);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h2, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0010__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0010__2 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0010__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module131;
    method Action rdReq_infoRam__0010__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__0010__1 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0010__1 ();
endinterface

module mkModule131 (Module131);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h1, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0010__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0010__1 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0010__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module132;
    method Action rdReq_infoRam__0010__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__0010__0 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0010__0 ();
endinterface

module mkModule132 (Module132);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h0, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0010__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0010__0 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0010__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module133;
    method Action rdReq_dataRam__0010 (Bit#(10) x_0);
    method Action wrReq_dataRam__0010 (Struct73 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0010 ();
endinterface

module mkModule133 (Module133);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__0010 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__0010 (Struct73 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0010 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module134;
    method Action rdReq_repRam__0010 (Bit#(8) x_0);
    method Action wrReq_repRam__0010 (Struct76 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0010 ();
endinterface

module mkModule134 (Module134);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h0, 8'h0, 8'h0, 8'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__0010 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__0010 (Struct76 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0010 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module135;
    method ActionValue#(Struct63) getMSHR_0010 (Bit#(3) x_0);
    method ActionValue#(Struct57) getPRqSlot_0010 (Struct56 x_0);
    method ActionValue#(Struct57) getCRqSlot_0010 (Struct56 x_0);
    method ActionValue#(Struct58) getWait_0010 ();
    method Action registerUL_0010 (Struct65 x_0);
    method Action registerDL_0010 (Struct77 x_0);
    method ActionValue#(Bit#(3)) getULImm_0010 (Struct1 x_0);
    method ActionValue#(Bit#(3)) getULCount_0010 ();
    method Action transferUpDown_0010 (Struct78 x_0);
    method ActionValue#(Bit#(3)) findUL_0010 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) findDL_0010 (Bit#(64) x_0);
    method Action releaseMSHR_0010 (Bit#(3) x_0);
    method Action addRs_0010 (Struct6 x_0);
    method ActionValue#(Struct59) getRsReady_0010 ();
endinterface

module mkModule135
    (Module135);
    Reg#(Vector#(6, Struct63)) rqs_0010 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct63) getMSHR_0010 (Bit#(3) x_0);
        let x_1 = (rqs_0010);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct57) getPRqSlot_0010 (Struct56 x_0);
        let x_1 = (rqs_0010);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0010 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct57) getCRqSlot_0010 (Struct56 x_0);
        let x_1 = (rqs_0010);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0010 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct58) getWait_0010 ();
        let x_1 = (rqs_0010);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        let x_6 = ?;
        if ((x_2).valid) begin
            Bit#(3) x_3 = ((x_2).data);
            Struct63 x_4 = ((x_1)[x_3]);
            rqs_0010 <= update (x_1, x_3, Struct63 {m_status :
            (Bit#(2))'(2'h3), m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul,
            m_msg : (x_4).m_msg, m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb,
            m_dl_rss_from : (x_4).m_dl_rss_from, m_dl_rss_recv :
            (x_4).m_dl_rss_recv, m_dl_rss : (x_4).m_dl_rss});
            Struct56 x_5 = (Struct56 {r_id : x_3, r_msg : (x_4).m_msg,
            r_msg_from : (x_4).m_qidx});
            x_6 = Struct58 {valid : (Bool)'(True), data : x_5};
        end else begin
            x_6 = Struct58 {valid : (Bool)'(False), data : unpack(0)};
        end
        return x_6;
    endmethod

    method Action registerUL_0010 (Struct65 x_0);
        let x_1 = (rqs_0010);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_0010 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_0010 (Struct77 x_0);
        let x_1 = (rqs_0010);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0010 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) getULImm_0010 (Struct1 x_0);
        let x_1 = (rqs_0010);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h6)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h7)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        rqs_0010 <= update (x_1, x_3, Struct63 {m_status : (Bit#(2))'(2'h3),
        m_next : Struct10 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul
        : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0), m_rsb :
        (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
        m_dl_rss : unpack(0)});
        return x_3;
    endmethod

    method ActionValue#(Bit#(3)) getULCount_0010 ();
        let x_1 = (rqs_0010);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h3)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + (((((x_1)[(Bit#(3))'(3'h4)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h5)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + ((Bit#(3))'(3'h0))))));
        return x_2;
    endmethod

    method Action transferUpDown_0010 (Struct78 x_0);
        let x_1 = (rqs_0010);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0010 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) findUL_0010 (Bit#(64) x_0);
        let x_1 = (rqs_0010);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))));
        return x_2;
    endmethod

    method ActionValue#(Bit#(3)) findDL_0010 (Bit#(64) x_0);
        let x_1 = (rqs_0010);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        return x_2;
    endmethod

    method Action releaseMSHR_0010 (Bit#(3) x_0);
        let x_1 = (rqs_0010);
        Struct63 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct63) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct63 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct63) x_6 = (update (x_3, x_4, Struct63 {m_status
            : (Bit#(2))'(2'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_0010 <= x_7;
    endmethod

    method Action addRs_0010 (Struct6 x_0);
        let x_1 = (rqs_0010);
        Bit#(64) x_2 = (((x_0).r_dl_msg).addr);
        Bit#(3) x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        Struct63 x_4 = ((x_1)[x_3]);
        Struct63 x_5 = (Struct63 {m_status : (x_4).m_status, m_next :
        (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg, m_qidx :
        (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : ((x_4).m_dl_rss_recv) |
        (((Bit#(2))'(2'h1)) << ((x_0).r_dl_midx)), m_dl_rss : update
        ((x_4).m_dl_rss, (x_0).r_dl_midx, (x_0).r_dl_msg)});
        rqs_0010 <= update (x_1, x_3, x_5);
    endmethod

    method ActionValue#(Struct59) getRsReady_0010 ();
        let x_1 = (rqs_0010);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h0)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h1)) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h2)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h3)) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h4)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h5)) :
        (unpack(0))))))))))))));
        Struct63 x_3 = ((x_1)[x_2]);
        Struct59 x_4 = (Struct59 {r_id : x_2, r_addr :
        ((x_3).m_msg).addr});
        return x_4;
    endmethod
endmodule

interface Module136;
    method Action enq_fifoInput0011 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoInput0011 ();
endinterface

module mkModule136 (Module136);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoInput0011 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoInput0011 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module137;
    method Action enq_fifoI2L0011 (Struct55 x_0);
    method ActionValue#(Struct55) deq_fifoI2L0011 ();
endinterface

module mkModule137 (Module137);
    FIFOF#(Struct55) pff <- mkFIFOF();

    method Action enq_fifoI2L0011 (Struct55 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct55) deq_fifoI2L0011 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module138;
    method Action enq_fifoL2E0011 (Struct62 x_0);
    method ActionValue#(Struct62) deq_fifoL2E0011 ();
endinterface

module mkModule138 (Module138);
    FIFOF#(Struct62) pff <- mkFIFOF();

    method Action enq_fifoL2E0011 (Struct62 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct62) deq_fifoL2E0011 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module139;
    method Action enq_fifo00110 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00110 ();
endinterface

module mkModule139 (Module139);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00110 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00110 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module140;
    method Action enq_fifo00111 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00111 ();
endinterface

module mkModule140 (Module140);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00111 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00111 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module141;
    method Action enq_fifo00112 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo00112 ();
endinterface

module mkModule141 (Module141);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo00112 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo00112 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module142;
    method Action enq_fifo001100 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo001100 ();
endinterface

module mkModule142 (Module142);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo001100 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo001100 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module143;
    method Action enq_fifo001102 (Struct1 x_0);
    method ActionValue#(Struct1) deq_fifo001102 ();
endinterface

module mkModule143 (Module143);
    FIFOF#(Struct1) pff <- mkFIFOF();

    method Action enq_fifo001102 (Struct1 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct1) deq_fifo001102 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module144;
    method Action enq_cp_1__0011 (Struct68 x_0);
    method ActionValue#(Struct68) deq_cp_1__0011 ();
endinterface

module mkModule144 (Module144);
    FIFOF#(Struct68) pff <- mkPipelineFIFOF();

    method Action enq_cp_1__0011 (Struct68 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct68) deq_cp_1__0011 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module145;
    method Action enq_cp_2__0011 (Struct69 x_0);
    method ActionValue#(Struct69) deq_cp_2__0011 ();
endinterface

module mkModule145 (Module145);
    FIFOF#(Struct69) pff <- mkPipelineFIFOF();

    method Action enq_cp_2__0011 (Struct69 x_0);
        pff.enq(x_0);
    endmethod

    method ActionValue#(Struct69) deq_cp_2__0011 ();
        pff.deq();
        return pff.first();
    endmethod

endmodule

interface Module146;
    method Action rdReq_infoRam__0011__3 (Bit#(8) x_0);
    method Action wrReq_infoRam__0011__3 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0011__3 ();
endinterface

module mkModule146 (Module146);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h3, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0011__3 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0011__3 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0011__3 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module147;
    method Action rdReq_infoRam__0011__2 (Bit#(8) x_0);
    method Action wrReq_infoRam__0011__2 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0011__2 ();
endinterface

module mkModule147 (Module147);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h2, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0011__2 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0011__2 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0011__2 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module148;
    method Action rdReq_infoRam__0011__1 (Bit#(8) x_0);
    method Action wrReq_infoRam__0011__1 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0011__1 ();
endinterface

module mkModule148 (Module148);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h1, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0011__1 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0011__1 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0011__1 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module149;
    method Action rdReq_infoRam__0011__0 (Bit#(8) x_0);
    method Action wrReq_infoRam__0011__0 (Struct72 x_0);
    method ActionValue#(Struct70) rdResp_infoRam__0011__0 ();
endinterface

module mkModule149 (Module149);
    RWBramCore#(Bit#(8), Struct70) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = Struct70 {tag: 51'h0, value: Struct11 {mesi_owned: False, mesi_status: 3'h1, mesi_dir_st: 3'h1, mesi_dir_sharers: 2'h0}};
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_infoRam__0011__0 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_infoRam__0011__0 (Struct72 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Struct70) rdResp_infoRam__0011__0 () if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module150;
    method Action rdReq_dataRam__0011 (Bit#(10) x_0);
    method Action wrReq_dataRam__0011 (Struct73 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0011 ();
endinterface

module mkModule150 (Module150);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(10)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(64'h0, 64'h0, 64'h0, 64'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_dataRam__0011 (Bit#(10) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_dataRam__0011 (Struct73 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0011 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module151;
    method Action rdReq_repRam__0011 (Bit#(8) x_0);
    method Action wrReq_repRam__0011 (Struct76 x_0);
    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0011 ();
endinterface

module mkModule151 (Module151);
    RWBramCore#(Bit#(8), Vector#(4, Bit#(8))) bram <- mkRWBramCore();
    Reg#(Bool) initDone <- mkReg(False);
    Reg#(Bit#(8)) initIdx <- mkReg(0);

    rule init (!initDone);
        let initData = vec(8'h0, 8'h0, 8'h0, 8'h0);
        bram.wrReq(initIdx, initData);
        initIdx <= initIdx + 1;
        initDone <= (initIdx == maxBound);
    endrule

    method Action rdReq_repRam__0011 (Bit#(8) x_0) if(initDone);
        bram.rdReq(x_0);
    endmethod

    method Action wrReq_repRam__0011 (Struct76 x_0) if(initDone);
        bram.wrReq(x_0.addr, x_0.datain);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0011 ()
    if(initDone);
        bram.deqRdResp ();
        let data = bram.rdResp ();
        return data;
    endmethod


endmodule

interface Module152;
    method ActionValue#(Struct63) getMSHR_0011 (Bit#(3) x_0);
    method ActionValue#(Struct57) getPRqSlot_0011 (Struct56 x_0);
    method ActionValue#(Struct57) getCRqSlot_0011 (Struct56 x_0);
    method ActionValue#(Struct58) getWait_0011 ();
    method Action registerUL_0011 (Struct65 x_0);
    method Action registerDL_0011 (Struct77 x_0);
    method ActionValue#(Bit#(3)) getULImm_0011 (Struct1 x_0);
    method ActionValue#(Bit#(3)) getULCount_0011 ();
    method Action transferUpDown_0011 (Struct78 x_0);
    method ActionValue#(Bit#(3)) findUL_0011 (Bit#(64) x_0);
    method ActionValue#(Bit#(3)) findDL_0011 (Bit#(64) x_0);
    method Action releaseMSHR_0011 (Bit#(3) x_0);
    method Action addRs_0011 (Struct6 x_0);
    method ActionValue#(Struct59) getRsReady_0011 ();
endinterface

module mkModule152
    (Module152);
    Reg#(Vector#(6, Struct63)) rqs_0011 <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Struct63) getMSHR_0011 (Bit#(3) x_0);
        let x_1 = (rqs_0011);
        return (x_1)[x_0];
    endmethod

    method ActionValue#(Struct57) getPRqSlot_0011 (Struct56 x_0);
        let x_1 = (rqs_0011);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0011 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct57) getCRqSlot_0011 (Struct56 x_0);
        let x_1 = (rqs_0011);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        Bool x_3 = ((x_2).valid);
        Bit#(3) x_4 = ((x_2).data);
        Bit#(64) x_5 = (((x_0).r_msg).addr);
        Struct10 x_6 = ((((! ((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h0)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h0)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h1)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h1)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h2)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h2)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h3)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h3)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h4)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h4)}) : ((((!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h0)))) && (!
        ((((x_1)[(Bit#(3))'(3'h5)]).m_next).valid))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_5)) ? (Struct10
        {valid : (Bool)'(True), data : (Bit#(3))'(3'h5)}) : (Struct10 {valid
        : (Bool)'(False), data : unpack(0)})))))))))))));
        Bool x_7 = ((x_6).valid);
        Bit#(3) x_8 = ((x_6).data);
        Struct57 x_9 = (Struct57 {s_has_slot : x_3, s_conflict : x_7, s_id :
        x_4});
        if (x_3) begin
            Struct63 x_10 = ((x_1)[x_8]);
            rqs_0011 <= update (update (x_1, x_4, Struct63 {m_status : (x_7 ?
            ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h3))), m_next : Struct10
            {valid : (Bool)'(False), data : unpack(0)}, m_is_ul : unpack(0),
            m_msg : (x_0).r_msg, m_qidx : (x_0).r_msg_from, m_rsb :
            unpack(0), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
            m_dl_rss : unpack(0)}), x_8, Struct63 {m_status :
            (x_10).m_status, m_next : (x_7 ? (Struct10 {valid :
            (Bool)'(True), data : x_4}) : ((x_10).m_next)), m_is_ul :
            (x_10).m_is_ul, m_msg : (x_10).m_msg, m_qidx : (x_10).m_qidx,
            m_rsb : (x_10).m_rsb, m_dl_rss_from : (x_10).m_dl_rss_from,
            m_dl_rss_recv : (x_10).m_dl_rss_recv, m_dl_rss :
            (x_10).m_dl_rss});
        end else begin

        end
        return x_9;
    endmethod

    method ActionValue#(Struct58) getWait_0011 ();
        let x_1 = (rqs_0011);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h0)}) : (((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h1)}) : (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h2)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h3)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h2)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))))))));
        let x_6 = ?;
        if ((x_2).valid) begin
            Bit#(3) x_3 = ((x_2).data);
            Struct63 x_4 = ((x_1)[x_3]);
            rqs_0011 <= update (x_1, x_3, Struct63 {m_status :
            (Bit#(2))'(2'h3), m_next : (x_4).m_next, m_is_ul : (x_4).m_is_ul,
            m_msg : (x_4).m_msg, m_qidx : (x_4).m_qidx, m_rsb : (x_4).m_rsb,
            m_dl_rss_from : (x_4).m_dl_rss_from, m_dl_rss_recv :
            (x_4).m_dl_rss_recv, m_dl_rss : (x_4).m_dl_rss});
            Struct56 x_5 = (Struct56 {r_id : x_3, r_msg : (x_4).m_msg,
            r_msg_from : (x_4).m_qidx});
            x_6 = Struct58 {valid : (Bool)'(True), data : x_5};
        end else begin
            x_6 = Struct58 {valid : (Bool)'(False), data : unpack(0)};
        end
        return x_6;
    endmethod

    method Action registerUL_0011 (Struct65 x_0);
        let x_1 = (rqs_0011);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(True), m_msg : (x_3).m_msg, m_qidx :
        zeroExtend((x_0).r_ul_rsbTo), m_rsb : (x_0).r_ul_rsb, m_dl_rss_from :
        unpack(0), m_dl_rss_recv : unpack(0), m_dl_rss : unpack(0)});
        rqs_0011 <= update (x_1, x_2, x_4);
    endmethod

    method Action registerDL_0011 (Struct77 x_0);
        let x_1 = (rqs_0011);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_0).r_dl_rsbTo, m_rsb : (x_0).r_dl_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0011 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) getULImm_0011 (Struct1 x_0);
        let x_1 = (rqs_0011);
        Struct10 x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h4)}) : (((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h5)}) : (((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h6)}) : (((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h0)) ? (Struct10 {valid : (Bool)'(True), data :
        (Bit#(3))'(3'h7)}) : (Struct10 {valid : (Bool)'(False), data :
        unpack(0)})))))))));
        when ((x_2).valid, noAction);
        Bit#(3) x_3 = ((x_2).data);
        rqs_0011 <= update (x_1, x_3, Struct63 {m_status : (Bit#(2))'(2'h3),
        m_next : Struct10 {valid : (Bool)'(False), data : unpack(0)}, m_is_ul
        : (Bool)'(True), m_msg : x_0, m_qidx : unpack(0), m_rsb :
        (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv : unpack(0),
        m_dl_rss : unpack(0)});
        return x_3;
    endmethod

    method ActionValue#(Bit#(3)) getULCount_0011 ();
        let x_1 = (rqs_0011);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h2)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h3)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + (((((x_1)[(Bit#(3))'(3'h4)]).m_is_ul ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((x_1)[(Bit#(3))'(3'h5)]).m_is_ul ? ((Bit#(3))'(3'h1)) :
        ((Bit#(3))'(3'h0)))) + ((Bit#(3))'(3'h0))))));
        return x_2;
    endmethod

    method Action transferUpDown_0011 (Struct78 x_0);
        let x_1 = (rqs_0011);
        Bit#(3) x_2 = ((x_0).r_id);
        Struct63 x_3 = ((x_1)[x_2]);
        Struct63 x_4 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        (x_3).m_next, m_is_ul : (Bool)'(False), m_msg : (x_3).m_msg, m_qidx :
        (x_3).m_qidx, m_rsb : (x_3).m_rsb, m_dl_rss_from :
        (x_0).r_dl_rss_from, m_dl_rss_recv : unpack(0), m_dl_rss :
        unpack(0)});
        rqs_0011 <= update (x_1, x_2, x_4);
    endmethod

    method ActionValue#(Bit#(3)) findUL_0011 (Bit#(64) x_0);
        let x_1 = (rqs_0011);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul)) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))));
        return x_2;
    endmethod

    method ActionValue#(Bit#(3)) findDL_0011 (Bit#(64) x_0);
        let x_1 = (rqs_0011);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        return x_2;
    endmethod

    method Action releaseMSHR_0011 (Bit#(3) x_0);
        let x_1 = (rqs_0011);
        Struct63 x_2 = ((x_1)[x_0]);
        Vector#(6, Struct63) x_3 = (update (x_1, x_0,
        unpack(0)));
        let x_7 = ?;
        if (((x_2).m_next).valid) begin
            Bit#(3) x_4 = (((x_2).m_next).data);
            Struct63 x_5 = ((x_1)[x_4]);
            Vector#(6, Struct63) x_6 = (update (x_3, x_4, Struct63 {m_status
            : (Bit#(2))'(2'h2), m_next : (x_5).m_next, m_is_ul :
            (x_5).m_is_ul, m_msg : (x_5).m_msg, m_qidx : (x_5).m_qidx, m_rsb
            : (x_5).m_rsb, m_dl_rss_from : (x_5).m_dl_rss_from, m_dl_rss_recv
            : (x_5).m_dl_rss_recv, m_dl_rss : (x_5).m_dl_rss}));
            x_7 = x_6;
        end else begin
            x_7 = x_3;
        end
        rqs_0011 <= x_7;
    endmethod

    method Action addRs_0011 (Struct6 x_0);
        let x_1 = (rqs_0011);
        Bit#(64) x_2 = (((x_0).r_dl_msg).addr);
        Bit#(3) x_3 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h0)) : (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h1)) : (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h2)) : (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h3)) : (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h4)) : (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).m_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h5)) : (unpack(0))))))))))))));
        Struct63 x_4 = ((x_1)[x_3]);
        Struct63 x_5 = (Struct63 {m_status : (x_4).m_status, m_next :
        (x_4).m_next, m_is_ul : (x_4).m_is_ul, m_msg : (x_4).m_msg, m_qidx :
        (x_4).m_qidx, m_rsb : (x_4).m_rsb, m_dl_rss_from :
        (x_4).m_dl_rss_from, m_dl_rss_recv : ((x_4).m_dl_rss_recv) |
        (((Bit#(2))'(2'h1)) << ((x_0).r_dl_midx)), m_dl_rss : update
        ((x_4).m_dl_rss, (x_0).r_dl_midx, (x_0).r_dl_msg)});
        rqs_0011 <= update (x_1, x_3, x_5);
    endmethod

    method ActionValue#(Struct59) getRsReady_0011 ();
        let x_1 = (rqs_0011);
        Bit#(3) x_2 = (((((((x_1)[(Bit#(3))'(3'h0)]).m_status) ==
        ((Bit#(2))'(2'h3))) && (! (((x_1)[(Bit#(3))'(3'h0)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h0)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h0)) :
        (((((((x_1)[(Bit#(3))'(3'h1)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h1)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h1)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h1)) :
        (((((((x_1)[(Bit#(3))'(3'h2)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h2)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h2)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h2)) :
        (((((((x_1)[(Bit#(3))'(3'h3)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h3)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h3)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h3)) :
        (((((((x_1)[(Bit#(3))'(3'h4)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h4)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h4)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h4)) :
        (((((((x_1)[(Bit#(3))'(3'h5)]).m_status) == ((Bit#(2))'(2'h3))) && (!
        (((x_1)[(Bit#(3))'(3'h5)]).m_is_ul))) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_from) ==
        (((x_1)[(Bit#(3))'(3'h5)]).m_dl_rss_recv)) ? ((Bit#(3))'(3'h5)) :
        (unpack(0))))))))))))));
        Struct63 x_3 = ((x_1)[x_2]);
        Struct59 x_4 = (Struct59 {r_id : x_2, r_addr :
        ((x_3).m_msg).addr});
        return x_4;
    endmethod
endmodule

interface Module153;

endinterface

module mkModule153#(function ActionValue#(Struct1) deq_fifo0010(),
    function Action enq_fifoCRqInput00(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0000())
    (Module153);
    Reg#(Bit#(1)) rr_00 <- mkReg(unpack(0));

    rule inc_rr_00;
        let x_0 = (rr_00);
        rr_00 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_00;
        let x_0 = (rr_00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo0000();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h0), ch_msg : x_1});
        let x_3 <- enq_fifoCRqInput00(x_2);
    endrule

    rule accept1_00;
        let x_0 = (rr_00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo0010();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h1), ch_msg : x_1});
        let x_3 <- enq_fifoCRqInput00(x_2);
    endrule

    // No methods in this module
endmodule

interface Module154;

endinterface

module mkModule154#(function ActionValue#(Struct1) deq_fifo0010(),
    function Action enq_fifoCRsInput00(Struct2 _),
    function ActionValue#(Struct1) deq_fifo0000())
    (Module154);
    Reg#(Bit#(1)) rr_00 <- mkReg(unpack(0));

    rule inc_rr_00;
        let x_0 = (rr_00);
        rr_00 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_00;
        let x_0 = (rr_00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo0000();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h0), ch_msg : x_1});
        let x_3 <- enq_fifoCRsInput00(x_2);
    endrule

    rule accept1_00;
        let x_0 = (rr_00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo0010();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h1), ch_msg : x_1});
        let x_3 <- enq_fifoCRsInput00(x_2);
    endrule

    // No methods in this module
endmodule

interface Module155;

endinterface

module mkModule155#(function ActionValue#(Struct2) deq_fifoCRsInput00(),
    function ActionValue#(Struct2) deq_fifoCRqInput00(),
    function Action enq_fifoInput00(Struct3 _),
    function ActionValue#(Struct1) deq_fifo002())
    (Module155);
    Reg#(Bit#(2)) rr_00 <- mkReg(unpack(0));

    rule inc_rr_00;
        let x_0 = (rr_00);
        rr_00 <= ((x_0) == ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h0)) : ((x_0) +
        ((Bit#(2))'(2'h1))));
    endrule

    rule accept0_00;
        let x_0 = (rr_00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 <- deq_fifo002();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg : x_1,
        ir_msg_from : {((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}, ir_mshr_id :
        unpack(0)});
        let x_3 <- enq_fifoInput00(x_2);
    endrule

    rule accept1_00;
        let x_0 = (rr_00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 <- deq_fifoCRqInput00();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_1).ch_msg, ir_msg_from : {((Bit#(2))'(2'h0)),((x_1).ch_idx)},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput00(x_2);
    endrule

    rule accept2_00;
        let x_0 = (rr_00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 <- deq_fifoCRsInput00();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_1).ch_msg, ir_msg_from : {((Bit#(2))'(2'h1)),((x_1).ch_idx)},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput00(x_2);
    endrule

    // No methods in this module
endmodule

interface Module156;
    method Action makeEnq_parentChildren00 (Struct17 x_0);
    method Action broadcast_parentChildren00 (Struct20 x_0);
endinterface

module mkModule156#(function Action enq_fifo0002(Struct1 _),
    function Action enq_fifo0012(Struct1 _),
    function Action enq_fifo001(Struct1 _),
    function Action enq_fifo000(Struct1 _))
    (Module156);

    // No rules in this module

    method Action makeEnq_parentChildren00 (Struct17 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo000((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo001((x_0).enq_msg);
            end else begin
                Bit#(1) x_3 = ((x_0).enq_ch_idx);
                Struct1 x_4 =
                ((x_0).enq_msg);
                if ((x_3) == ((Bit#(1))'(1'h1))) begin
                    let x_5 <- enq_fifo0012(x_4);
                end else
                    begin
                    if ((x_3) == ((Bit#(1))'(1'h0))) begin
                        let x_6 <- enq_fifo0002(x_4);
                    end else begin

                    end
                end
            end
        end
    endmethod

    method Action broadcast_parentChildren00 (Struct20 x_0);
        Bit#(2) x_1 = ((x_0).cs_inds);
        Struct1 x_2 =
        ((x_0).cs_msg);
        if (((x_1) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == (x_1))
            begin
            let x_3 <- enq_fifo0012(x_2);
        end else begin

        end
        if (((x_1) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == (x_1))
            begin
            let x_5 <- enq_fifo0002(x_2);
        end else begin

        end
    endmethod
endmodule

interface Module157;
    method Action repGetRq__00 (Bit#(10) x_0);
    method ActionValue#(Vector#(16, Bit#(8))) repGetRs__00 ();
    method Action repAccess__00 (Struct35 x_0);
endinterface

module mkModule157#(function Action wrReq_repRam__00(Struct39 _),
    function ActionValue#(Vector#(16, Bit#(8))) rdResp_repRam__00(),
    function Action rdReq_repRam__00(Bit#(10) _))
    (Module157);

    // No rules in this module

    method Action repGetRq__00 (Bit#(10) x_0);
        let x_1 <- rdReq_repRam__00(x_0);
    endmethod

    method ActionValue#(Vector#(16, Bit#(8))) repGetRs__00 ();
        let x_1 <- rdResp_repRam__00();
        return x_1;
    endmethod

    method Action repAccess__00 (Struct35 x_0);
        Vector#(16, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(4))'(4'hf)]) +
        (((((x_1)[(Bit#(4))'(4'hf)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(4))'(4'hf)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_3 = (update (x_1, (Bit#(4))'(4'hf),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(4))'(4'he)]) +
        (((((x_3)[(Bit#(4))'(4'he)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(4))'(4'he)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_5 = (update (x_3, (Bit#(4))'(4'he),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(4))'(4'hd)]) +
        (((((x_5)[(Bit#(4))'(4'hd)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(4))'(4'hd)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_7 = (update (x_5, (Bit#(4))'(4'hd),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(4))'(4'hc)]) +
        (((((x_7)[(Bit#(4))'(4'hc)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(4))'(4'hc)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_9 = (update (x_7, (Bit#(4))'(4'hc),
        x_8));
        Bit#(8) x_10 = (((x_9)[(Bit#(4))'(4'hb)]) +
        (((((x_9)[(Bit#(4))'(4'hb)]) == ((Bit#(8))'(8'h0))) ||
        (((x_9)[(Bit#(4))'(4'hb)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_11 = (update (x_9, (Bit#(4))'(4'hb),
        x_10));
        Bit#(8) x_12 = (((x_11)[(Bit#(4))'(4'ha)]) +
        (((((x_11)[(Bit#(4))'(4'ha)]) == ((Bit#(8))'(8'h0))) ||
        (((x_11)[(Bit#(4))'(4'ha)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_13 = (update (x_11, (Bit#(4))'(4'ha),
        x_12));
        Bit#(8) x_14 = (((x_13)[(Bit#(4))'(4'h9)]) +
        (((((x_13)[(Bit#(4))'(4'h9)]) == ((Bit#(8))'(8'h0))) ||
        (((x_13)[(Bit#(4))'(4'h9)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_15 = (update (x_13, (Bit#(4))'(4'h9),
        x_14));
        Bit#(8) x_16 = (((x_15)[(Bit#(4))'(4'h8)]) +
        (((((x_15)[(Bit#(4))'(4'h8)]) == ((Bit#(8))'(8'h0))) ||
        (((x_15)[(Bit#(4))'(4'h8)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_17 = (update (x_15, (Bit#(4))'(4'h8),
        x_16));
        Bit#(8) x_18 = (((x_17)[(Bit#(4))'(4'h7)]) +
        (((((x_17)[(Bit#(4))'(4'h7)]) == ((Bit#(8))'(8'h0))) ||
        (((x_17)[(Bit#(4))'(4'h7)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_19 = (update (x_17, (Bit#(4))'(4'h7),
        x_18));
        Bit#(8) x_20 = (((x_19)[(Bit#(4))'(4'h6)]) +
        (((((x_19)[(Bit#(4))'(4'h6)]) == ((Bit#(8))'(8'h0))) ||
        (((x_19)[(Bit#(4))'(4'h6)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_21 = (update (x_19, (Bit#(4))'(4'h6),
        x_20));
        Bit#(8) x_22 = (((x_21)[(Bit#(4))'(4'h5)]) +
        (((((x_21)[(Bit#(4))'(4'h5)]) == ((Bit#(8))'(8'h0))) ||
        (((x_21)[(Bit#(4))'(4'h5)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_23 = (update (x_21, (Bit#(4))'(4'h5),
        x_22));
        Bit#(8) x_24 = (((x_23)[(Bit#(4))'(4'h4)]) +
        (((((x_23)[(Bit#(4))'(4'h4)]) == ((Bit#(8))'(8'h0))) ||
        (((x_23)[(Bit#(4))'(4'h4)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_25 = (update (x_23, (Bit#(4))'(4'h4),
        x_24));
        Bit#(8) x_26 = (((x_25)[(Bit#(4))'(4'h3)]) +
        (((((x_25)[(Bit#(4))'(4'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_25)[(Bit#(4))'(4'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_27 = (update (x_25, (Bit#(4))'(4'h3),
        x_26));
        Bit#(8) x_28 = (((x_27)[(Bit#(4))'(4'h2)]) +
        (((((x_27)[(Bit#(4))'(4'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_27)[(Bit#(4))'(4'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_29 = (update (x_27, (Bit#(4))'(4'h2),
        x_28));
        Bit#(8) x_30 = (((x_29)[(Bit#(4))'(4'h1)]) +
        (((((x_29)[(Bit#(4))'(4'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_29)[(Bit#(4))'(4'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_31 = (update (x_29, (Bit#(4))'(4'h1),
        x_30));
        Bit#(8) x_32 = (((x_31)[(Bit#(4))'(4'h0)]) +
        (((((x_31)[(Bit#(4))'(4'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_31)[(Bit#(4))'(4'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(16, Bit#(8)) x_33 = (update (x_31, (Bit#(4))'(4'h0),
        x_32));
        let x_36 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(16, Bit#(8)) x_34 = (update (x_33, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_36 = x_34;
        end else begin
            Vector#(16, Bit#(8)) x_35 = (update (x_33, (x_0).acc_way,
            (Bit#(8))'(8'hff)));
            x_36 = x_35;
        end
        Struct39 x_37 = (Struct39 {addr : (x_0).acc_index, datain :
        x_36});
        let x_38 <- wrReq_repRam__00(x_37);
    endmethod
endmodule

interface Module158;

endinterface

module mkModule158#(function ActionValue#(Struct1) deq_fifo00010(),
    function Action enq_fifoCRqInput000(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00000())
    (Module158);
    Reg#(Bit#(1)) rr_000 <- mkReg(unpack(0));

    rule inc_rr_000;
        let x_0 = (rr_000);
        rr_000 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_000;
        let x_0 = (rr_000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00000();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h0), ch_msg : x_1});
        let x_3 <- enq_fifoCRqInput000(x_2);
    endrule

    rule accept1_000;
        let x_0 = (rr_000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo00010();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h1), ch_msg : x_1});
        let x_3 <- enq_fifoCRqInput000(x_2);
    endrule

    // No methods in this module
endmodule

interface Module159;

endinterface

module mkModule159#(function ActionValue#(Struct1) deq_fifo00010(),
    function Action enq_fifoCRsInput000(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00000())
    (Module159);
    Reg#(Bit#(1)) rr_000 <- mkReg(unpack(0));

    rule inc_rr_000;
        let x_0 = (rr_000);
        rr_000 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_000;
        let x_0 = (rr_000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00000();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h0), ch_msg : x_1});
        let x_3 <- enq_fifoCRsInput000(x_2);
    endrule

    rule accept1_000;
        let x_0 = (rr_000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo00010();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h1), ch_msg : x_1});
        let x_3 <- enq_fifoCRsInput000(x_2);
    endrule

    // No methods in this module
endmodule

interface Module160;

endinterface

module mkModule160#(function ActionValue#(Struct2) deq_fifoCRsInput000(),
    function ActionValue#(Struct2) deq_fifoCRqInput000(),
    function Action enq_fifoInput000(Struct3 _),
    function ActionValue#(Struct1) deq_fifo0002())
    (Module160);
    Reg#(Bit#(2)) rr_000 <- mkReg(unpack(0));

    rule inc_rr_000;
        let x_0 = (rr_000);
        rr_000 <= ((x_0) == ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h0)) : ((x_0)
        + ((Bit#(2))'(2'h1))));
    endrule

    rule accept0_000;
        let x_0 = (rr_000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 <- deq_fifo0002();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg : x_1,
        ir_msg_from : {((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}, ir_mshr_id :
        unpack(0)});
        let x_3 <- enq_fifoInput000(x_2);
    endrule

    rule accept1_000;
        let x_0 = (rr_000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 <- deq_fifoCRqInput000();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_1).ch_msg, ir_msg_from : {((Bit#(2))'(2'h0)),((x_1).ch_idx)},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput000(x_2);
    endrule

    rule accept2_000;
        let x_0 = (rr_000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 <- deq_fifoCRsInput000();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_1).ch_msg, ir_msg_from : {((Bit#(2))'(2'h1)),((x_1).ch_idx)},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput000(x_2);
    endrule

    // No methods in this module
endmodule

interface Module161;
    method Action makeEnq_parentChildren000 (Struct17 x_0);
    method Action broadcast_parentChildren000 (Struct20 x_0);
endinterface

module mkModule161#(function Action enq_fifo00002(Struct1 _),
    function Action enq_fifo00012(Struct1 _),
    function Action enq_fifo0001(Struct1 _),
    function Action enq_fifo0000(Struct1 _))
    (Module161);

    // No rules in this module

    method Action makeEnq_parentChildren000 (Struct17 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo0000((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo0001((x_0).enq_msg);
            end else begin
                Bit#(1) x_3 = ((x_0).enq_ch_idx);
                Struct1 x_4 =
                ((x_0).enq_msg);
                if ((x_3) == ((Bit#(1))'(1'h1))) begin
                    let x_5 <- enq_fifo00012(x_4);
                end else
                    begin
                    if ((x_3) == ((Bit#(1))'(1'h0))) begin
                        let x_6 <- enq_fifo00002(x_4);
                    end else begin

                    end
                end
            end
        end
    endmethod

    method Action broadcast_parentChildren000 (Struct20 x_0);
        Bit#(2) x_1 = ((x_0).cs_inds);
        Struct1 x_2 =
        ((x_0).cs_msg);
        if (((x_1) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == (x_1))
            begin
            let x_3 <- enq_fifo00012(x_2);
        end else begin

        end
        if (((x_1) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == (x_1))
            begin
            let x_5 <- enq_fifo00002(x_2);
        end else begin

        end
    endmethod
endmodule

interface Module162;
    method Action repGetRq__000 (Bit#(9) x_0);
    method ActionValue#(Vector#(8, Bit#(8))) repGetRs__000 ();
    method Action repAccess__000 (Struct51 x_0);
endinterface

module mkModule162#(function Action wrReq_repRam__000(Struct54 _),
    function ActionValue#(Vector#(8, Bit#(8))) rdResp_repRam__000(),
    function Action rdReq_repRam__000(Bit#(9) _))
    (Module162);

    // No rules in this module

    method Action repGetRq__000 (Bit#(9) x_0);
        let x_1 <- rdReq_repRam__000(x_0);
    endmethod

    method ActionValue#(Vector#(8, Bit#(8))) repGetRs__000 ();
        let x_1 <- rdResp_repRam__000();
        return x_1;
    endmethod

    method Action repAccess__000 (Struct51 x_0);
        Vector#(8, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(3))'(3'h7)]) +
        (((((x_1)[(Bit#(3))'(3'h7)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(3))'(3'h7)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_3 = (update (x_1, (Bit#(3))'(3'h7),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(3))'(3'h6)]) +
        (((((x_3)[(Bit#(3))'(3'h6)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(3))'(3'h6)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_5 = (update (x_3, (Bit#(3))'(3'h6),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(3))'(3'h5)]) +
        (((((x_5)[(Bit#(3))'(3'h5)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(3))'(3'h5)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_7 = (update (x_5, (Bit#(3))'(3'h5),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(3))'(3'h4)]) +
        (((((x_7)[(Bit#(3))'(3'h4)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(3))'(3'h4)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_9 = (update (x_7, (Bit#(3))'(3'h4),
        x_8));
        Bit#(8) x_10 = (((x_9)[(Bit#(3))'(3'h3)]) +
        (((((x_9)[(Bit#(3))'(3'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_9)[(Bit#(3))'(3'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_11 = (update (x_9, (Bit#(3))'(3'h3),
        x_10));
        Bit#(8) x_12 = (((x_11)[(Bit#(3))'(3'h2)]) +
        (((((x_11)[(Bit#(3))'(3'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_11)[(Bit#(3))'(3'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_13 = (update (x_11, (Bit#(3))'(3'h2),
        x_12));
        Bit#(8) x_14 = (((x_13)[(Bit#(3))'(3'h1)]) +
        (((((x_13)[(Bit#(3))'(3'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_13)[(Bit#(3))'(3'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_15 = (update (x_13, (Bit#(3))'(3'h1),
        x_14));
        Bit#(8) x_16 = (((x_15)[(Bit#(3))'(3'h0)]) +
        (((((x_15)[(Bit#(3))'(3'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_15)[(Bit#(3))'(3'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_17 = (update (x_15, (Bit#(3))'(3'h0),
        x_16));
        let x_20 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(8, Bit#(8)) x_18 = (update (x_17, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_20 = x_18;
        end else begin
            Vector#(8, Bit#(8)) x_19 = (update (x_17, (x_0).acc_way,
            (Bit#(8))'(8'hff)));
            x_20 = x_19;
        end
        Struct54 x_21 = (Struct54 {addr : (x_0).acc_index, datain :
        x_20});
        let x_22 <- wrReq_repRam__000(x_21);
    endmethod
endmodule

interface Module163;

endinterface

module mkModule163#(function ActionValue#(Struct1) deq_fifo000000(),
    function Action enq_fifoInput0000(Struct55 _),
    function ActionValue#(Struct1) deq_fifo00002())
    (Module163);
    Reg#(Bit#(1)) rr_0000 <- mkReg(unpack(0));

    rule inc_rr_0000;
        let x_0 = (rr_0000);
        rr_0000 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_0000;
        let x_0 = (rr_0000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00002();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0000(x_2);
    endrule

    rule accept1_0000;
        let x_0 = (rr_0000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo000000();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h0)),((Bit#(1))'(1'h0))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0000(x_2);
    endrule

    // No methods in this module
endmodule

interface Module164;
    method Action makeEnq_parentChildren0000 (Struct17 x_0);
endinterface

module mkModule164#(function Action enq_fifo000002(Struct1 _),
    function Action enq_fifo00001(Struct1 _),
    function Action enq_fifo00000(Struct1 _))
    (Module164);

    // No rules in this module

    method Action makeEnq_parentChildren0000 (Struct17 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo00000((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo00001((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo000002(x_3);
            end
        end
    endmethod
endmodule

interface Module165;
    method Action repGetRq__0000 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0000 ();
    method Action repAccess__0000 (Struct74 x_0);
endinterface

module mkModule165#(function Action wrReq_repRam__0000(Struct76 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0000(),
    function Action rdReq_repRam__0000(Bit#(8) _))
    (Module165);

    // No rules in this module

    method Action repGetRq__0000 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__0000(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0000 ();
        let x_1 <- rdResp_repRam__0000();
        return x_1;
    endmethod

    method Action repAccess__0000 (Struct74 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'hff)));
            x_12 = x_11;
        end
        Struct76 x_13 = (Struct76 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__0000(x_13);
    endmethod
endmodule

interface Module166;

endinterface

module mkModule166#(function ActionValue#(Struct1) deq_fifo000100(),
    function Action enq_fifoInput0001(Struct55 _),
    function ActionValue#(Struct1) deq_fifo00012())
    (Module166);
    Reg#(Bit#(1)) rr_0001 <- mkReg(unpack(0));

    rule inc_rr_0001;
        let x_0 = (rr_0001);
        rr_0001 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_0001;
        let x_0 = (rr_0001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00012();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0001(x_2);
    endrule

    rule accept1_0001;
        let x_0 = (rr_0001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo000100();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h0)),((Bit#(1))'(1'h0))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0001(x_2);
    endrule

    // No methods in this module
endmodule

interface Module167;
    method Action makeEnq_parentChildren0001 (Struct17 x_0);
endinterface

module mkModule167#(function Action enq_fifo000102(Struct1 _),
    function Action enq_fifo00011(Struct1 _),
    function Action enq_fifo00010(Struct1 _))
    (Module167);

    // No rules in this module

    method Action makeEnq_parentChildren0001 (Struct17 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo00010((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo00011((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo000102(x_3);
            end
        end
    endmethod
endmodule

interface Module168;
    method Action repGetRq__0001 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0001 ();
    method Action repAccess__0001 (Struct74 x_0);
endinterface

module mkModule168#(function Action wrReq_repRam__0001(Struct76 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0001(),
    function Action rdReq_repRam__0001(Bit#(8) _))
    (Module168);

    // No rules in this module

    method Action repGetRq__0001 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__0001(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0001 ();
        let x_1 <- rdResp_repRam__0001();
        return x_1;
    endmethod

    method Action repAccess__0001 (Struct74 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'hff)));
            x_12 = x_11;
        end
        Struct76 x_13 = (Struct76 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__0001(x_13);
    endmethod
endmodule

interface Module169;

endinterface

module mkModule169#(function ActionValue#(Struct1) deq_fifo00110(),
    function Action enq_fifoCRqInput001(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00100())
    (Module169);
    Reg#(Bit#(1)) rr_001 <- mkReg(unpack(0));

    rule inc_rr_001;
        let x_0 = (rr_001);
        rr_001 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_001;
        let x_0 = (rr_001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00100();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h0), ch_msg : x_1});
        let x_3 <- enq_fifoCRqInput001(x_2);
    endrule

    rule accept1_001;
        let x_0 = (rr_001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo00110();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h1), ch_msg : x_1});
        let x_3 <- enq_fifoCRqInput001(x_2);
    endrule

    // No methods in this module
endmodule

interface Module170;

endinterface

module mkModule170#(function ActionValue#(Struct1) deq_fifo00110(),
    function Action enq_fifoCRsInput001(Struct2 _),
    function ActionValue#(Struct1) deq_fifo00100())
    (Module170);
    Reg#(Bit#(1)) rr_001 <- mkReg(unpack(0));

    rule inc_rr_001;
        let x_0 = (rr_001);
        rr_001 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_001;
        let x_0 = (rr_001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00100();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h0), ch_msg : x_1});
        let x_3 <- enq_fifoCRsInput001(x_2);
    endrule

    rule accept1_001;
        let x_0 = (rr_001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo00110();
        Struct2 x_2 = (Struct2 {ch_idx : (Bit#(1))'(1'h1), ch_msg : x_1});
        let x_3 <- enq_fifoCRsInput001(x_2);
    endrule

    // No methods in this module
endmodule

interface Module171;

endinterface

module mkModule171#(function ActionValue#(Struct2) deq_fifoCRsInput001(),
    function ActionValue#(Struct2) deq_fifoCRqInput001(),
    function Action enq_fifoInput001(Struct3 _),
    function ActionValue#(Struct1) deq_fifo0012())
    (Module171);
    Reg#(Bit#(2)) rr_001 <- mkReg(unpack(0));

    rule inc_rr_001;
        let x_0 = (rr_001);
        rr_001 <= ((x_0) == ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h0)) : ((x_0)
        + ((Bit#(2))'(2'h1))));
    endrule

    rule accept0_001;
        let x_0 = (rr_001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 <- deq_fifo0012();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg : x_1,
        ir_msg_from : {((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}, ir_mshr_id :
        unpack(0)});
        let x_3 <- enq_fifoInput001(x_2);
    endrule

    rule accept1_001;
        let x_0 = (rr_001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 <- deq_fifoCRqInput001();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_1).ch_msg, ir_msg_from : {((Bit#(2))'(2'h0)),((x_1).ch_idx)},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput001(x_2);
    endrule

    rule accept2_001;
        let x_0 = (rr_001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 <- deq_fifoCRsInput001();
        Struct3 x_2 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_1).ch_msg, ir_msg_from : {((Bit#(2))'(2'h1)),((x_1).ch_idx)},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput001(x_2);
    endrule

    // No methods in this module
endmodule

interface Module172;
    method Action makeEnq_parentChildren001 (Struct17 x_0);
    method Action broadcast_parentChildren001 (Struct20 x_0);
endinterface

module mkModule172#(function Action enq_fifo00102(Struct1 _),
    function Action enq_fifo00112(Struct1 _),
    function Action enq_fifo0011(Struct1 _),
    function Action enq_fifo0010(Struct1 _))
    (Module172);

    // No rules in this module

    method Action makeEnq_parentChildren001 (Struct17 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo0010((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo0011((x_0).enq_msg);
            end else begin
                Bit#(1) x_3 = ((x_0).enq_ch_idx);
                Struct1 x_4 =
                ((x_0).enq_msg);
                if ((x_3) == ((Bit#(1))'(1'h1))) begin
                    let x_5 <- enq_fifo00112(x_4);
                end else
                    begin
                    if ((x_3) == ((Bit#(1))'(1'h0))) begin
                        let x_6 <- enq_fifo00102(x_4);
                    end else begin

                    end
                end
            end
        end
    endmethod

    method Action broadcast_parentChildren001 (Struct20 x_0);
        Bit#(2) x_1 = ((x_0).cs_inds);
        Struct1 x_2 =
        ((x_0).cs_msg);
        if (((x_1) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == (x_1))
            begin
            let x_3 <- enq_fifo00112(x_2);
        end else begin

        end
        if (((x_1) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == (x_1))
            begin
            let x_5 <- enq_fifo00102(x_2);
        end else begin

        end
    endmethod
endmodule

interface Module173;
    method Action repGetRq__001 (Bit#(9) x_0);
    method ActionValue#(Vector#(8, Bit#(8))) repGetRs__001 ();
    method Action repAccess__001 (Struct51 x_0);
endinterface

module mkModule173#(function Action wrReq_repRam__001(Struct54 _),
    function ActionValue#(Vector#(8, Bit#(8))) rdResp_repRam__001(),
    function Action rdReq_repRam__001(Bit#(9) _))
    (Module173);

    // No rules in this module

    method Action repGetRq__001 (Bit#(9) x_0);
        let x_1 <- rdReq_repRam__001(x_0);
    endmethod

    method ActionValue#(Vector#(8, Bit#(8))) repGetRs__001 ();
        let x_1 <- rdResp_repRam__001();
        return x_1;
    endmethod

    method Action repAccess__001 (Struct51 x_0);
        Vector#(8, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(3))'(3'h7)]) +
        (((((x_1)[(Bit#(3))'(3'h7)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(3))'(3'h7)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_3 = (update (x_1, (Bit#(3))'(3'h7),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(3))'(3'h6)]) +
        (((((x_3)[(Bit#(3))'(3'h6)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(3))'(3'h6)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_5 = (update (x_3, (Bit#(3))'(3'h6),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(3))'(3'h5)]) +
        (((((x_5)[(Bit#(3))'(3'h5)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(3))'(3'h5)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_7 = (update (x_5, (Bit#(3))'(3'h5),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(3))'(3'h4)]) +
        (((((x_7)[(Bit#(3))'(3'h4)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(3))'(3'h4)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_9 = (update (x_7, (Bit#(3))'(3'h4),
        x_8));
        Bit#(8) x_10 = (((x_9)[(Bit#(3))'(3'h3)]) +
        (((((x_9)[(Bit#(3))'(3'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_9)[(Bit#(3))'(3'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_11 = (update (x_9, (Bit#(3))'(3'h3),
        x_10));
        Bit#(8) x_12 = (((x_11)[(Bit#(3))'(3'h2)]) +
        (((((x_11)[(Bit#(3))'(3'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_11)[(Bit#(3))'(3'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_13 = (update (x_11, (Bit#(3))'(3'h2),
        x_12));
        Bit#(8) x_14 = (((x_13)[(Bit#(3))'(3'h1)]) +
        (((((x_13)[(Bit#(3))'(3'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_13)[(Bit#(3))'(3'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_15 = (update (x_13, (Bit#(3))'(3'h1),
        x_14));
        Bit#(8) x_16 = (((x_15)[(Bit#(3))'(3'h0)]) +
        (((((x_15)[(Bit#(3))'(3'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_15)[(Bit#(3))'(3'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(8, Bit#(8)) x_17 = (update (x_15, (Bit#(3))'(3'h0),
        x_16));
        let x_20 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(8, Bit#(8)) x_18 = (update (x_17, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_20 = x_18;
        end else begin
            Vector#(8, Bit#(8)) x_19 = (update (x_17, (x_0).acc_way,
            (Bit#(8))'(8'hff)));
            x_20 = x_19;
        end
        Struct54 x_21 = (Struct54 {addr : (x_0).acc_index, datain :
        x_20});
        let x_22 <- wrReq_repRam__001(x_21);
    endmethod
endmodule

interface Module174;

endinterface

module mkModule174#(function ActionValue#(Struct1) deq_fifo001000(),
    function Action enq_fifoInput0010(Struct55 _),
    function ActionValue#(Struct1) deq_fifo00102())
    (Module174);
    Reg#(Bit#(1)) rr_0010 <- mkReg(unpack(0));

    rule inc_rr_0010;
        let x_0 = (rr_0010);
        rr_0010 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_0010;
        let x_0 = (rr_0010);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00102();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0010(x_2);
    endrule

    rule accept1_0010;
        let x_0 = (rr_0010);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo001000();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h0)),((Bit#(1))'(1'h0))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0010(x_2);
    endrule

    // No methods in this module
endmodule

interface Module175;
    method Action makeEnq_parentChildren0010 (Struct17 x_0);
endinterface

module mkModule175#(function Action enq_fifo001002(Struct1 _),
    function Action enq_fifo00101(Struct1 _),
    function Action enq_fifo00100(Struct1 _))
    (Module175);

    // No rules in this module

    method Action makeEnq_parentChildren0010 (Struct17 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo00100((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo00101((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo001002(x_3);
            end
        end
    endmethod
endmodule

interface Module176;
    method Action repGetRq__0010 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0010 ();
    method Action repAccess__0010 (Struct74 x_0);
endinterface

module mkModule176#(function Action wrReq_repRam__0010(Struct76 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0010(),
    function Action rdReq_repRam__0010(Bit#(8) _))
    (Module176);

    // No rules in this module

    method Action repGetRq__0010 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__0010(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0010 ();
        let x_1 <- rdResp_repRam__0010();
        return x_1;
    endmethod

    method Action repAccess__0010 (Struct74 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'hff)));
            x_12 = x_11;
        end
        Struct76 x_13 = (Struct76 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__0010(x_13);
    endmethod
endmodule

interface Module177;

endinterface

module mkModule177#(function ActionValue#(Struct1) deq_fifo001100(),
    function Action enq_fifoInput0011(Struct55 _),
    function ActionValue#(Struct1) deq_fifo00112())
    (Module177);
    Reg#(Bit#(1)) rr_0011 <- mkReg(unpack(0));

    rule inc_rr_0011;
        let x_0 = (rr_0011);
        rr_0011 <= (x_0) + ((Bit#(1))'(1'h1));
    endrule

    rule accept0_0011;
        let x_0 = (rr_0011);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 <- deq_fifo00112();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0011(x_2);
    endrule

    rule accept1_0011;
        let x_0 = (rr_0011);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 <- deq_fifo001100();
        Struct55 x_2 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_1, ir_msg_from : {((Bit#(2))'(2'h0)),((Bit#(1))'(1'h0))},
        ir_mshr_id : unpack(0)});
        let x_3 <- enq_fifoInput0011(x_2);
    endrule

    // No methods in this module
endmodule

interface Module178;
    method Action makeEnq_parentChildren0011 (Struct17 x_0);
endinterface

module mkModule178#(function Action enq_fifo001102(Struct1 _),
    function Action enq_fifo00111(Struct1 _),
    function Action enq_fifo00110(Struct1 _))
    (Module178);

    // No rules in this module

    method Action makeEnq_parentChildren0011 (Struct17 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
            let x_1 <- enq_fifo00110((x_0).enq_msg);
        end else
            begin
            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
                let x_2 <- enq_fifo00111((x_0).enq_msg);
            end else begin
                Struct1 x_3 = ((x_0).enq_msg);
                let x_4 <- enq_fifo001102(x_3);
            end
        end
    endmethod
endmodule

interface Module179;
    method Action repGetRq__0011 (Bit#(8) x_0);
    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0011 ();
    method Action repAccess__0011 (Struct74 x_0);
endinterface

module mkModule179#(function Action wrReq_repRam__0011(Struct76 _),
    function ActionValue#(Vector#(4, Bit#(8))) rdResp_repRam__0011(),
    function Action rdReq_repRam__0011(Bit#(8) _))
    (Module179);

    // No rules in this module

    method Action repGetRq__0011 (Bit#(8) x_0);
        let x_1 <- rdReq_repRam__0011(x_0);
    endmethod

    method ActionValue#(Vector#(4, Bit#(8))) repGetRs__0011 ();
        let x_1 <- rdResp_repRam__0011();
        return x_1;
    endmethod

    method Action repAccess__0011 (Struct74 x_0);
        Vector#(4, Bit#(8)) x_1 = ((x_0).acc_reps);
        Bit#(8) x_2 = (((x_1)[(Bit#(2))'(2'h3)]) +
        (((((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'h0))) ||
        (((x_1)[(Bit#(2))'(2'h3)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_3 = (update (x_1, (Bit#(2))'(2'h3),
        x_2));
        Bit#(8) x_4 = (((x_3)[(Bit#(2))'(2'h2)]) +
        (((((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'h0))) ||
        (((x_3)[(Bit#(2))'(2'h2)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_5 = (update (x_3, (Bit#(2))'(2'h2),
        x_4));
        Bit#(8) x_6 = (((x_5)[(Bit#(2))'(2'h1)]) +
        (((((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'h0))) ||
        (((x_5)[(Bit#(2))'(2'h1)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_7 = (update (x_5, (Bit#(2))'(2'h1),
        x_6));
        Bit#(8) x_8 = (((x_7)[(Bit#(2))'(2'h0)]) +
        (((((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'h0))) ||
        (((x_7)[(Bit#(2))'(2'h0)]) == ((Bit#(8))'(8'hff))) ?
        ((Bit#(8))'(8'h0)) : ((Bit#(8))'(8'h1)))));
        Vector#(4, Bit#(8)) x_9 = (update (x_7, (Bit#(2))'(2'h0),
        x_8));
        let x_12 = ?;
        if (((x_0).acc_type) == ((Bit#(1))'(1'h0))) begin
            Vector#(4, Bit#(8)) x_10 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'h1)));
            x_12 = x_10;
        end else begin
            Vector#(4, Bit#(8)) x_11 = (update (x_9, (x_0).acc_way,
            (Bit#(8))'(8'hff)));
            x_12 = x_11;
        end
        Struct76 x_13 = (Struct76 {addr : (x_0).acc_index, datain :
        x_12});
        let x_14 <- wrReq_repRam__0011(x_13);
    endmethod
endmodule

interface Module180;
    method Action cache__00__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct9) cache__00__infoRsValueRq ();
    method ActionValue#(Vector#(4, Bit#(64))) cache__00__valueRsLineRq
    (Struct16 x_0);
    method ActionValue#(Struct23) cache__00__getVictim ();
    method Action cache__00__setVictimRq (Struct24 x_0);
    method ActionValue#(Bit#(4)) cache__00__releaseVictim (Bit#(64) x_0);
    method ActionValue#(Bit#(1)) cache__00__getVictimCount ();
endinterface

module mkModule180#(function Action wrReq_edirRam__00__7(Struct37 _),
    function Action wrReq_edirRam__00__6(Struct37 _),
    function Action wrReq_edirRam__00__5(Struct37 _),
    function Action wrReq_edirRam__00__4(Struct37 _),
    function Action wrReq_edirRam__00__3(Struct37 _),
    function Action wrReq_edirRam__00__2(Struct37 _),
    function Action wrReq_edirRam__00__1(Struct37 _),
    function Action wrReq_edirRam__00__0(Struct37 _),
    function Action wrReq_dataRam__00(Struct36 _),
    function Action repAccess__00(Struct35 _),
    function Action wrReq_infoRam__00__15(Struct34 _),
    function Action wrReq_infoRam__00__14(Struct34 _),
    function Action wrReq_infoRam__00__13(Struct34 _),
    function Action wrReq_infoRam__00__12(Struct34 _),
    function Action wrReq_infoRam__00__11(Struct34 _),
    function Action wrReq_infoRam__00__10(Struct34 _),
    function Action wrReq_infoRam__00__9(Struct34 _),
    function Action wrReq_infoRam__00__8(Struct34 _),
    function Action wrReq_infoRam__00__7(Struct34 _),
    function Action wrReq_infoRam__00__6(Struct34 _),
    function Action wrReq_infoRam__00__5(Struct34 _),
    function Action wrReq_infoRam__00__4(Struct34 _),
    function Action wrReq_infoRam__00__3(Struct34 _),
    function Action wrReq_infoRam__00__2(Struct34 _),
    function Action wrReq_infoRam__00__1(Struct34 _),
    function Action wrReq_infoRam__00__0(Struct34 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__00(),
    function ActionValue#(Struct27) deq_cp_2__00(),
    function Action rdReq_dataRam__00(Bit#(14) _),
    function ActionValue#(Vector#(16, Bit#(8))) repGetRs__00(),
    function ActionValue#(Struct31) rdResp_edirRam__00__7(),
    function ActionValue#(Struct31) rdResp_edirRam__00__6(),
    function ActionValue#(Struct31) rdResp_edirRam__00__5(),
    function ActionValue#(Struct31) rdResp_edirRam__00__4(),
    function ActionValue#(Struct31) rdResp_edirRam__00__3(),
    function ActionValue#(Struct31) rdResp_edirRam__00__2(),
    function ActionValue#(Struct31) rdResp_edirRam__00__1(),
    function ActionValue#(Struct31) rdResp_edirRam__00__0(),
    function ActionValue#(Struct29) rdResp_infoRam__00__15(),
    function ActionValue#(Struct29) rdResp_infoRam__00__14(),
    function ActionValue#(Struct29) rdResp_infoRam__00__13(),
    function ActionValue#(Struct29) rdResp_infoRam__00__12(),
    function ActionValue#(Struct29) rdResp_infoRam__00__11(),
    function ActionValue#(Struct29) rdResp_infoRam__00__10(),
    function ActionValue#(Struct29) rdResp_infoRam__00__9(),
    function ActionValue#(Struct29) rdResp_infoRam__00__8(),
    function ActionValue#(Struct29) rdResp_infoRam__00__7(),
    function ActionValue#(Struct29) rdResp_infoRam__00__6(),
    function ActionValue#(Struct29) rdResp_infoRam__00__5(),
    function ActionValue#(Struct29) rdResp_infoRam__00__4(),
    function ActionValue#(Struct29) rdResp_infoRam__00__3(),
    function ActionValue#(Struct29) rdResp_infoRam__00__2(),
    function ActionValue#(Struct29) rdResp_infoRam__00__1(),
    function ActionValue#(Struct29) rdResp_infoRam__00__0(),
    function Action enq_cp_2__00(Struct27 _),
    function ActionValue#(Struct25) deq_cp_1__00(),
    function Action repGetRq__00(Bit#(10) _),
    function Action rdReq_edirRam__00__7(Bit#(10) _),
    function Action rdReq_edirRam__00__6(Bit#(10) _),
    function Action rdReq_edirRam__00__5(Bit#(10) _),
    function Action rdReq_edirRam__00__4(Bit#(10) _),
    function Action rdReq_edirRam__00__3(Bit#(10) _),
    function Action rdReq_edirRam__00__2(Bit#(10) _),
    function Action rdReq_edirRam__00__1(Bit#(10) _),
    function Action rdReq_edirRam__00__0(Bit#(10) _),
    function Action rdReq_infoRam__00__15(Bit#(10) _),
    function Action rdReq_infoRam__00__14(Bit#(10) _),
    function Action rdReq_infoRam__00__13(Bit#(10) _),
    function Action rdReq_infoRam__00__12(Bit#(10) _),
    function Action rdReq_infoRam__00__11(Bit#(10) _),
    function Action rdReq_infoRam__00__10(Bit#(10) _),
    function Action rdReq_infoRam__00__9(Bit#(10) _),
    function Action rdReq_infoRam__00__8(Bit#(10) _),
    function Action rdReq_infoRam__00__7(Bit#(10) _),
    function Action rdReq_infoRam__00__6(Bit#(10) _),
    function Action rdReq_infoRam__00__5(Bit#(10) _),
    function Action rdReq_infoRam__00__4(Bit#(10) _),
    function Action rdReq_infoRam__00__3(Bit#(10) _),
    function Action rdReq_infoRam__00__2(Bit#(10) _),
    function Action rdReq_infoRam__00__1(Bit#(10) _),
    function Action rdReq_infoRam__00__0(Bit#(10) _),
    function Action enq_cp_1__00(Struct25 _))
    (Module180);
    Reg#(Vector#(4, Struct23)) victims__00 <- mkReg(unpack(0));

    // No rules in this module

    method Action cache__00__infoRq (Bit#(64) x_0);
        let x_1 = (victims__00);
        Struct23 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            let x_3 <- enq_cp_1__00(Struct25 {tag : (x_0)[63:15], index :
            (x_0)[14:5], victim_found : Struct26 {valid : (Bool)'(True), data
            : (Bit#(1))'(1'h0)}});
        end else begin
            Struct23 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                let x_5 <- enq_cp_1__00(Struct25 {tag : (x_0)[63:15], index :
                (x_0)[14:5], victim_found : Struct26 {valid : (Bool)'(True),
                data : (Bit#(1))'(1'h1)}});
            end else begin
                Struct23 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    let x_7 <- enq_cp_1__00(Struct25 {tag : (x_0)[63:15],
                    index : (x_0)[14:5], victim_found : Struct26 {valid :
                    (Bool)'(True), data : (Bit#(1))'(1'h0)}});
                end else begin
                    Struct23 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        let x_9 <- enq_cp_1__00(Struct25 {tag : (x_0)[63:15],
                        index : (x_0)[14:5], victim_found : Struct26 {valid :
                        (Bool)'(True), data : (Bit#(1))'(1'h1)}});
                    end else begin
                        Bit#(10) x_10 = ((x_0)[14:5]);
                        let x_11 <- rdReq_infoRam__00__0(x_10);
                        let x_12 <- rdReq_infoRam__00__1(x_10);
                        let x_13 <- rdReq_infoRam__00__2(x_10);
                        let x_14 <- rdReq_infoRam__00__3(x_10);
                        let x_15 <- rdReq_infoRam__00__4(x_10);
                        let x_16 <- rdReq_infoRam__00__5(x_10);
                        let x_17 <- rdReq_infoRam__00__6(x_10);
                        let x_18 <- rdReq_infoRam__00__7(x_10);
                        let x_19 <- rdReq_infoRam__00__8(x_10);
                        let x_20 <- rdReq_infoRam__00__9(x_10);
                        let x_21 <- rdReq_infoRam__00__10(x_10);
                        let x_22 <- rdReq_infoRam__00__11(x_10);
                        let x_23 <- rdReq_infoRam__00__12(x_10);
                        let x_24 <- rdReq_infoRam__00__13(x_10);
                        let x_25 <- rdReq_infoRam__00__14(x_10);
                        let x_26 <- rdReq_infoRam__00__15(x_10);
                        let x_27 <- rdReq_edirRam__00__0(x_10);
                        let x_28 <- rdReq_edirRam__00__1(x_10);
                        let x_29 <- rdReq_edirRam__00__2(x_10);
                        let x_30 <- rdReq_edirRam__00__3(x_10);
                        let x_31 <- rdReq_edirRam__00__4(x_10);
                        let x_32 <- rdReq_edirRam__00__5(x_10);
                        let x_33 <- rdReq_edirRam__00__6(x_10);
                        let x_34 <- rdReq_edirRam__00__7(x_10);
                        let x_35 <- repGetRq__00(x_10);
                        let x_36 <- enq_cp_1__00(Struct25 {tag :
                        (x_0)[63:15], index : (x_0)[14:5], victim_found :
                        Struct26 {valid : (Bool)'(False), data :
                        unpack(0)}});
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Struct9) cache__00__infoRsValueRq ();
        let x_1 <- deq_cp_1__00();
        Bit#(49) x_2 = ((x_1).tag);
        Bit#(10) x_3 =
        ((x_1).index);
        let x_104 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_4 = (((x_1).victim_found).data);
            let x_5 = (victims__00);
            Struct23 x_6 = ((x_5)[x_4]);
            Struct9 x_7 = (Struct9 {info_index : x_3, info_hit :
            (Bool)'(True), info_way : unpack(0), edir_hit : (Bool)'(False),
            edir_way : unpack(0), edir_slot : Struct10 {valid :
            (Bool)'(False), data : unpack(0)}, info : (x_6).victim_info});
            let x_8 <- enq_cp_2__00(Struct27 {victim_found :
            (x_1).victim_found, may_victim : unpack(0), reps :
            unpack(0)});
            x_104 = x_7;
        end else begin
            Vector#(16, Struct29) x_9 = (unpack(0));
            let x_10 <- rdResp_infoRam__00__0();
            Vector#(16, Struct29) x_11 = (update (x_9, (Bit#(4))'(4'h0),
            x_10));
            let x_12 <- rdResp_infoRam__00__1();
            Vector#(16, Struct29) x_13 = (update (x_11, (Bit#(4))'(4'h1),
            x_12));
            let x_14 <- rdResp_infoRam__00__2();
            Vector#(16, Struct29) x_15 = (update (x_13, (Bit#(4))'(4'h2),
            x_14));
            let x_16 <- rdResp_infoRam__00__3();
            Vector#(16, Struct29) x_17 = (update (x_15, (Bit#(4))'(4'h3),
            x_16));
            let x_18 <- rdResp_infoRam__00__4();
            Vector#(16, Struct29) x_19 = (update (x_17, (Bit#(4))'(4'h4),
            x_18));
            let x_20 <- rdResp_infoRam__00__5();
            Vector#(16, Struct29) x_21 = (update (x_19, (Bit#(4))'(4'h5),
            x_20));
            let x_22 <- rdResp_infoRam__00__6();
            Vector#(16, Struct29) x_23 = (update (x_21, (Bit#(4))'(4'h6),
            x_22));
            let x_24 <- rdResp_infoRam__00__7();
            Vector#(16, Struct29) x_25 = (update (x_23, (Bit#(4))'(4'h7),
            x_24));
            let x_26 <- rdResp_infoRam__00__8();
            Vector#(16, Struct29) x_27 = (update (x_25, (Bit#(4))'(4'h8),
            x_26));
            let x_28 <- rdResp_infoRam__00__9();
            Vector#(16, Struct29) x_29 = (update (x_27, (Bit#(4))'(4'h9),
            x_28));
            let x_30 <- rdResp_infoRam__00__10();
            Vector#(16, Struct29) x_31 = (update (x_29, (Bit#(4))'(4'ha),
            x_30));
            let x_32 <- rdResp_infoRam__00__11();
            Vector#(16, Struct29) x_33 = (update (x_31, (Bit#(4))'(4'hb),
            x_32));
            let x_34 <- rdResp_infoRam__00__12();
            Vector#(16, Struct29) x_35 = (update (x_33, (Bit#(4))'(4'hc),
            x_34));
            let x_36 <- rdResp_infoRam__00__13();
            Vector#(16, Struct29) x_37 = (update (x_35, (Bit#(4))'(4'hd),
            x_36));
            let x_38 <- rdResp_infoRam__00__14();
            Vector#(16, Struct29) x_39 = (update (x_37, (Bit#(4))'(4'he),
            x_38));
            let x_40 <- rdResp_infoRam__00__15();
            Vector#(16, Struct29) x_41 = (update (x_39, (Bit#(4))'(4'hf),
            x_40));
            Struct30 x_42 = (((((x_41)[(Bit#(4))'(4'h0)]).tag) == (x_2) ?
            (Struct30 {tm_hit : (Bool)'(True), tm_way : (Bit#(4))'(4'h0),
            tm_value : ((x_41)[(Bit#(4))'(4'h0)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h1)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h1), tm_value :
            ((x_41)[(Bit#(4))'(4'h1)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h2)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h2), tm_value :
            ((x_41)[(Bit#(4))'(4'h2)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h3)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h3), tm_value :
            ((x_41)[(Bit#(4))'(4'h3)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h4)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h4), tm_value :
            ((x_41)[(Bit#(4))'(4'h4)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h5)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h5), tm_value :
            ((x_41)[(Bit#(4))'(4'h5)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h6)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h6), tm_value :
            ((x_41)[(Bit#(4))'(4'h6)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h7)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h7), tm_value :
            ((x_41)[(Bit#(4))'(4'h7)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h8)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h8), tm_value :
            ((x_41)[(Bit#(4))'(4'h8)]).value}) :
            (((((x_41)[(Bit#(4))'(4'h9)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'h9), tm_value :
            ((x_41)[(Bit#(4))'(4'h9)]).value}) :
            (((((x_41)[(Bit#(4))'(4'ha)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'ha), tm_value :
            ((x_41)[(Bit#(4))'(4'ha)]).value}) :
            (((((x_41)[(Bit#(4))'(4'hb)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'hb), tm_value :
            ((x_41)[(Bit#(4))'(4'hb)]).value}) :
            (((((x_41)[(Bit#(4))'(4'hc)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'hc), tm_value :
            ((x_41)[(Bit#(4))'(4'hc)]).value}) :
            (((((x_41)[(Bit#(4))'(4'hd)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'hd), tm_value :
            ((x_41)[(Bit#(4))'(4'hd)]).value}) :
            (((((x_41)[(Bit#(4))'(4'he)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'he), tm_value :
            ((x_41)[(Bit#(4))'(4'he)]).value}) :
            (((((x_41)[(Bit#(4))'(4'hf)]).tag) == (x_2) ? (Struct30 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(4))'(4'hf), tm_value :
            ((x_41)[(Bit#(4))'(4'hf)]).value}) :
            (unpack(0))))))))))))))))))))))))))))))))));
            Vector#(8, Struct31) x_43 = (unpack(0));
            let x_44 <- rdResp_edirRam__00__0();
            Vector#(8, Struct31) x_45 = (update (x_43, (Bit#(3))'(3'h0),
            x_44));
            let x_46 <- rdResp_edirRam__00__1();
            Vector#(8, Struct31) x_47 = (update (x_45, (Bit#(3))'(3'h1),
            x_46));
            let x_48 <- rdResp_edirRam__00__2();
            Vector#(8, Struct31) x_49 = (update (x_47, (Bit#(3))'(3'h2),
            x_48));
            let x_50 <- rdResp_edirRam__00__3();
            Vector#(8, Struct31) x_51 = (update (x_49, (Bit#(3))'(3'h3),
            x_50));
            let x_52 <- rdResp_edirRam__00__4();
            Vector#(8, Struct31) x_53 = (update (x_51, (Bit#(3))'(3'h4),
            x_52));
            let x_54 <- rdResp_edirRam__00__5();
            Vector#(8, Struct31) x_55 = (update (x_53, (Bit#(3))'(3'h5),
            x_54));
            let x_56 <- rdResp_edirRam__00__6();
            Vector#(8, Struct31) x_57 = (update (x_55, (Bit#(3))'(3'h6),
            x_56));
            let x_58 <- rdResp_edirRam__00__7();
            Vector#(8, Struct31) x_59 = (update (x_57, (Bit#(3))'(3'h7),
            x_58));
            Struct33 x_60 = (((((x_59)[(Bit#(3))'(3'h0)]).tag) == (x_2) ?
            (Struct33 {tm_hit : (Bool)'(True), tm_way : (Bit#(3))'(3'h0),
            tm_value : ((x_59)[(Bit#(3))'(3'h0)]).value}) :
            (((((x_59)[(Bit#(3))'(3'h1)]).tag) == (x_2) ? (Struct33 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h1), tm_value :
            ((x_59)[(Bit#(3))'(3'h1)]).value}) :
            (((((x_59)[(Bit#(3))'(3'h2)]).tag) == (x_2) ? (Struct33 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h2), tm_value :
            ((x_59)[(Bit#(3))'(3'h2)]).value}) :
            (((((x_59)[(Bit#(3))'(3'h3)]).tag) == (x_2) ? (Struct33 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h3), tm_value :
            ((x_59)[(Bit#(3))'(3'h3)]).value}) :
            (((((x_59)[(Bit#(3))'(3'h4)]).tag) == (x_2) ? (Struct33 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h4), tm_value :
            ((x_59)[(Bit#(3))'(3'h4)]).value}) :
            (((((x_59)[(Bit#(3))'(3'h5)]).tag) == (x_2) ? (Struct33 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h5), tm_value :
            ((x_59)[(Bit#(3))'(3'h5)]).value}) :
            (((((x_59)[(Bit#(3))'(3'h6)]).tag) == (x_2) ? (Struct33 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h6), tm_value :
            ((x_59)[(Bit#(3))'(3'h6)]).value}) :
            (((((x_59)[(Bit#(3))'(3'h7)]).tag) == (x_2) ? (Struct33 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h7), tm_value :
            ((x_59)[(Bit#(3))'(3'h7)]).value}) :
            (unpack(0))))))))))))))))));
            Struct32 x_61 = ((x_60).tm_value);
            Struct10 x_62 =
            (((((((x_59)[(Bit#(3))'(3'h0)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h0)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h0)}) :
            (((((((x_59)[(Bit#(3))'(3'h1)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h1)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h1)}) :
            (((((((x_59)[(Bit#(3))'(3'h2)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h2)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h2)}) :
            (((((((x_59)[(Bit#(3))'(3'h3)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h3)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h3)}) :
            (((((((x_59)[(Bit#(3))'(3'h4)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h4)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h4)}) :
            (((((((x_59)[(Bit#(3))'(3'h5)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h5)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h5)}) :
            (((((((x_59)[(Bit#(3))'(3'h6)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h6)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h6)}) :
            (((((((x_59)[(Bit#(3))'(3'h7)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_59)[(Bit#(3))'(3'h7)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct10 {valid : (Bool)'(True), data :
            (Bit#(3))'(3'h7)}) : (Struct10 {valid : (Bool)'(False), data :
            unpack(0)})))))))))))))))));
            let x_63 <- repGetRs__00();
            Bit#(4) x_64 = (unpack(0));
            Bit#(8) x_65 = (unpack(0));
            Bit#(4) x_66 = ((! (((x_63)[(Bit#(4))'(4'hf)]) < (x_65)) ?
            ((Bit#(4))'(4'hf)) : (x_64)));
            Bit#(8) x_67 = ((! (((x_63)[(Bit#(4))'(4'hf)]) < (x_65)) ?
            ((x_63)[(Bit#(4))'(4'hf)]) : (x_65)));
            Bit#(4) x_68 = ((! (((x_63)[(Bit#(4))'(4'he)]) < (x_67)) ?
            ((Bit#(4))'(4'he)) : (x_66)));
            Bit#(8) x_69 = ((! (((x_63)[(Bit#(4))'(4'he)]) < (x_67)) ?
            ((x_63)[(Bit#(4))'(4'he)]) : (x_67)));
            Bit#(4) x_70 = ((! (((x_63)[(Bit#(4))'(4'hd)]) < (x_69)) ?
            ((Bit#(4))'(4'hd)) : (x_68)));
            Bit#(8) x_71 = ((! (((x_63)[(Bit#(4))'(4'hd)]) < (x_69)) ?
            ((x_63)[(Bit#(4))'(4'hd)]) : (x_69)));
            Bit#(4) x_72 = ((! (((x_63)[(Bit#(4))'(4'hc)]) < (x_71)) ?
            ((Bit#(4))'(4'hc)) : (x_70)));
            Bit#(8) x_73 = ((! (((x_63)[(Bit#(4))'(4'hc)]) < (x_71)) ?
            ((x_63)[(Bit#(4))'(4'hc)]) : (x_71)));
            Bit#(4) x_74 = ((! (((x_63)[(Bit#(4))'(4'hb)]) < (x_73)) ?
            ((Bit#(4))'(4'hb)) : (x_72)));
            Bit#(8) x_75 = ((! (((x_63)[(Bit#(4))'(4'hb)]) < (x_73)) ?
            ((x_63)[(Bit#(4))'(4'hb)]) : (x_73)));
            Bit#(4) x_76 = ((! (((x_63)[(Bit#(4))'(4'ha)]) < (x_75)) ?
            ((Bit#(4))'(4'ha)) : (x_74)));
            Bit#(8) x_77 = ((! (((x_63)[(Bit#(4))'(4'ha)]) < (x_75)) ?
            ((x_63)[(Bit#(4))'(4'ha)]) : (x_75)));
            Bit#(4) x_78 = ((! (((x_63)[(Bit#(4))'(4'h9)]) < (x_77)) ?
            ((Bit#(4))'(4'h9)) : (x_76)));
            Bit#(8) x_79 = ((! (((x_63)[(Bit#(4))'(4'h9)]) < (x_77)) ?
            ((x_63)[(Bit#(4))'(4'h9)]) : (x_77)));
            Bit#(4) x_80 = ((! (((x_63)[(Bit#(4))'(4'h8)]) < (x_79)) ?
            ((Bit#(4))'(4'h8)) : (x_78)));
            Bit#(8) x_81 = ((! (((x_63)[(Bit#(4))'(4'h8)]) < (x_79)) ?
            ((x_63)[(Bit#(4))'(4'h8)]) : (x_79)));
            Bit#(4) x_82 = ((! (((x_63)[(Bit#(4))'(4'h7)]) < (x_81)) ?
            ((Bit#(4))'(4'h7)) : (x_80)));
            Bit#(8) x_83 = ((! (((x_63)[(Bit#(4))'(4'h7)]) < (x_81)) ?
            ((x_63)[(Bit#(4))'(4'h7)]) : (x_81)));
            Bit#(4) x_84 = ((! (((x_63)[(Bit#(4))'(4'h6)]) < (x_83)) ?
            ((Bit#(4))'(4'h6)) : (x_82)));
            Bit#(8) x_85 = ((! (((x_63)[(Bit#(4))'(4'h6)]) < (x_83)) ?
            ((x_63)[(Bit#(4))'(4'h6)]) : (x_83)));
            Bit#(4) x_86 = ((! (((x_63)[(Bit#(4))'(4'h5)]) < (x_85)) ?
            ((Bit#(4))'(4'h5)) : (x_84)));
            Bit#(8) x_87 = ((! (((x_63)[(Bit#(4))'(4'h5)]) < (x_85)) ?
            ((x_63)[(Bit#(4))'(4'h5)]) : (x_85)));
            Bit#(4) x_88 = ((! (((x_63)[(Bit#(4))'(4'h4)]) < (x_87)) ?
            ((Bit#(4))'(4'h4)) : (x_86)));
            Bit#(8) x_89 = ((! (((x_63)[(Bit#(4))'(4'h4)]) < (x_87)) ?
            ((x_63)[(Bit#(4))'(4'h4)]) : (x_87)));
            Bit#(4) x_90 = ((! (((x_63)[(Bit#(4))'(4'h3)]) < (x_89)) ?
            ((Bit#(4))'(4'h3)) : (x_88)));
            Bit#(8) x_91 = ((! (((x_63)[(Bit#(4))'(4'h3)]) < (x_89)) ?
            ((x_63)[(Bit#(4))'(4'h3)]) : (x_89)));
            Bit#(4) x_92 = ((! (((x_63)[(Bit#(4))'(4'h2)]) < (x_91)) ?
            ((Bit#(4))'(4'h2)) : (x_90)));
            Bit#(8) x_93 = ((! (((x_63)[(Bit#(4))'(4'h2)]) < (x_91)) ?
            ((x_63)[(Bit#(4))'(4'h2)]) : (x_91)));
            Bit#(4) x_94 = ((! (((x_63)[(Bit#(4))'(4'h1)]) < (x_93)) ?
            ((Bit#(4))'(4'h1)) : (x_92)));
            Bit#(8) x_95 = ((! (((x_63)[(Bit#(4))'(4'h1)]) < (x_93)) ?
            ((x_63)[(Bit#(4))'(4'h1)]) : (x_93)));
            Bit#(4) x_96 = ((! (((x_63)[(Bit#(4))'(4'h0)]) < (x_95)) ?
            ((Bit#(4))'(4'h0)) : (x_94)));
            Bit#(8) x_97 = ((! (((x_63)[(Bit#(4))'(4'h0)]) < (x_95)) ?
            ((x_63)[(Bit#(4))'(4'h0)]) : (x_95)));
            Struct9 x_98 = (Struct9 {info_index : x_3, info_hit :
            (x_42).tm_hit, info_way : (x_42).tm_way, edir_hit :
            (x_60).tm_hit, edir_way : (x_60).tm_way, edir_slot : x_62, info :
            ((x_42).tm_hit ? ((x_42).tm_value) : (Struct11 {mesi_owned :
            (Bool)'(False), mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
            (x_61).mesi_edir_st, mesi_dir_sharers :
            (x_61).mesi_edir_sharers}))});
            Struct29 x_99 = ((x_41)[x_96]);
            Bit#(49) x_100 = ((x_99).tag);
            Struct11 x_101 = ((x_99).value);
            let x_102 <- enq_cp_2__00(Struct27 {victim_found : Struct26
            {valid : (Bool)'(False), data : unpack(0)}, may_victim : Struct28
            {mv_addr : {(x_100),({(x_3),((Bit#(5))'(5'h0))})}, mv_info :
            x_101}, reps : x_63});
            let x_103 <- rdReq_dataRam__00({(((x_42).tm_hit ? ((x_42).tm_way)
            : (x_96))),(x_3)});
            x_104 = x_98;
        end
        return x_104;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__00__valueRsLineRq
    (Struct16 x_0);
        let x_1 <- deq_cp_2__00();
        let x_2 =
        (victims__00);
        let x_93 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_3 = (((x_1).victim_found).data);
            Struct23 x_4 = ((x_2)[x_3]);
            Struct23 x_5 = (Struct23 {victim_valid : (Bool)'(True),
            victim_addr : (x_4).victim_addr, victim_info : ((x_0).info_write
            ? ((x_0).info) : ((x_4).victim_info)), victim_value :
            ((x_0).value_write ? ((x_0).value) : ((x_4).victim_value)),
            victim_req : (x_4).victim_req});
            victims__00 <= update (x_2, x_3, x_5);
            x_93 = (x_4).victim_value;
        end else begin
            let x_6 <- rdResp_dataRam__00();
            Bit#(64) x_7 = ((x_0).addr);
            Bit#(10) x_8 = ((x_7)[14:5]);
            Bit#(4) x_9 = ((x_0).info_way);
            Struct11 x_10 = ((x_0).info);
            Bool x_11 = ((! ((x_10).mesi_owned)) && (((x_10).mesi_status) ==
            ((Bit#(3))'(3'h1))));
            if ((((x_0).info_hit) || (! (x_11))) || ((! ((x_0).edir_hit)) &&
                (x_11)))
                begin
                if ((x_0).info_write) begin
                    Struct34 x_12 = (Struct34 {addr : x_8, datain : Struct29
                    {tag : (x_7)[63:15], value :
                    x_10}});
                    if ((x_9) == ((Bit#(4))'(4'h0))) begin
                        let x_13 <- wrReq_infoRam__00__0(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h1))) begin
                        let x_15 <- wrReq_infoRam__00__1(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h2))) begin
                        let x_17 <- wrReq_infoRam__00__2(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h3))) begin
                        let x_19 <- wrReq_infoRam__00__3(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h4))) begin
                        let x_21 <- wrReq_infoRam__00__4(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h5))) begin
                        let x_23 <- wrReq_infoRam__00__5(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h6))) begin
                        let x_25 <- wrReq_infoRam__00__6(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h7))) begin
                        let x_27 <- wrReq_infoRam__00__7(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h8))) begin
                        let x_29 <- wrReq_infoRam__00__8(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'h9))) begin
                        let x_31 <- wrReq_infoRam__00__9(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'ha))) begin
                        let x_33 <- wrReq_infoRam__00__10(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'hb))) begin
                        let x_35 <- wrReq_infoRam__00__11(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'hc))) begin
                        let x_37 <- wrReq_infoRam__00__12(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'hd))) begin
                        let x_39 <- wrReq_infoRam__00__13(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'he))) begin
                        let x_41 <- wrReq_infoRam__00__14(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(4))'(4'hf))) begin
                        let x_43 <- wrReq_infoRam__00__15(x_12);
                    end else begin

                    end
                    Struct28 x_45 = ((x_1).may_victim);
                    Struct26 x_46 = ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid
                    ? ((((x_2)[(Bit#(1))'(1'h0)]).victim_valid ?
                    ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid ? (Struct26
                    {valid : (Bool)'(False), data : unpack(0)}) : (Struct26
                    {valid : (Bool)'(True), data : (Bit#(1))'(1'h1)}))) :
                    (Struct26 {valid : (Bool)'(True), data :
                    (Bit#(1))'(1'h0)}))) : (Struct26 {valid : (Bool)'(True),
                    data : (Bit#(1))'(1'h1)})));
                    Bit#(1) x_47 = ((x_46).data);
                    victims__00 <= update (x_2, x_47, Struct23 {victim_valid
                    : (Bool)'(True), victim_addr : (x_45).mv_addr,
                    victim_info : (x_45).mv_info, victim_value : x_6,
                    victim_req : Struct14 {valid : (Bool)'(False), data :
                    unpack(0)}});
                    let x_48 <- repAccess__00(Struct35 {acc_type :
                    ((((x_10).mesi_dir_st) == ((Bit#(3))'(3'h0))) ||
                    (((x_10).mesi_dir_st) == ((Bit#(3))'(3'h1))) ?
                    ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))), acc_reps :
                    (x_1).reps, acc_index : x_8, acc_way : x_9});
                end else begin

                end
                if ((x_0).value_write) begin
                    Struct36 x_50 = (Struct36 {addr : {(x_9),((x_7)[14:5])},
                    datain : (x_0).value});
                    let x_51 <- wrReq_dataRam__00(x_50);
                end else begin

                end
            end else begin

            end
            if (((x_0).info_write) && ((x_0).edir_hit)) begin
                Bit#(3) x_54 = ((x_0).edir_way);
                Struct37 x_55 = (Struct37 {addr : (x_7)[14:5], datain :
                Struct31 {tag : (x_7)[63:15], value : (x_11 ? (Struct32
                {mesi_edir_st : (x_10).mesi_dir_st, mesi_edir_sharers :
                (x_10).mesi_dir_sharers}) :
                (unpack(0)))}});
                if ((x_54) == ((Bit#(3))'(3'h0))) begin
                    let x_56 <- wrReq_edirRam__00__0(x_55);
                end else begin

                end
                if ((x_54) == ((Bit#(3))'(3'h1))) begin
                    let x_58 <- wrReq_edirRam__00__1(x_55);
                end else begin

                end
                if ((x_54) == ((Bit#(3))'(3'h2))) begin
                    let x_60 <- wrReq_edirRam__00__2(x_55);
                end else begin

                end
                if ((x_54) == ((Bit#(3))'(3'h3))) begin
                    let x_62 <- wrReq_edirRam__00__3(x_55);
                end else begin

                end
                if ((x_54) == ((Bit#(3))'(3'h4))) begin
                    let x_64 <- wrReq_edirRam__00__4(x_55);
                end else begin

                end
                if ((x_54) == ((Bit#(3))'(3'h5))) begin
                    let x_66 <- wrReq_edirRam__00__5(x_55);
                end else begin

                end
                if ((x_54) == ((Bit#(3))'(3'h6))) begin
                    let x_68 <- wrReq_edirRam__00__6(x_55);
                end else begin

                end
                if ((x_54) == ((Bit#(3))'(3'h7))) begin
                    let x_70 <- wrReq_edirRam__00__7(x_55);
                end else begin

                end
            end else begin
                Struct10 x_72 =
                ((x_0).edir_slot);
                if (((! ((x_0).edir_hit)) && ((x_72).valid)) && (x_11))
                    begin
                    Bit#(3) x_73 = ((x_72).data);
                    Struct37 x_74 = (Struct37 {addr : (x_7)[14:5], datain :
                    Struct31 {tag : (x_7)[63:15], value : Struct32
                    {mesi_edir_st : (x_10).mesi_dir_st, mesi_edir_sharers :
                    (x_10).mesi_dir_sharers}}});
                    if ((x_73) == ((Bit#(3))'(3'h0))) begin
                        let x_75 <- wrReq_edirRam__00__0(x_74);
                    end else begin

                    end
                    if ((x_73) == ((Bit#(3))'(3'h1))) begin
                        let x_77 <- wrReq_edirRam__00__1(x_74);
                    end else begin

                    end
                    if ((x_73) == ((Bit#(3))'(3'h2))) begin
                        let x_79 <- wrReq_edirRam__00__2(x_74);
                    end else begin

                    end
                    if ((x_73) == ((Bit#(3))'(3'h3))) begin
                        let x_81 <- wrReq_edirRam__00__3(x_74);
                    end else begin

                    end
                    if ((x_73) == ((Bit#(3))'(3'h4))) begin
                        let x_83 <- wrReq_edirRam__00__4(x_74);
                    end else begin

                    end
                    if ((x_73) == ((Bit#(3))'(3'h5))) begin
                        let x_85 <- wrReq_edirRam__00__5(x_74);
                    end else begin

                    end
                    if ((x_73) == ((Bit#(3))'(3'h6))) begin
                        let x_87 <- wrReq_edirRam__00__6(x_74);
                    end else begin

                    end
                    if ((x_73) == ((Bit#(3))'(3'h7))) begin
                        let x_89 <- wrReq_edirRam__00__7(x_74);
                    end else begin

                    end
                end else begin

                end
            end
            x_93 = x_6;
        end
        return x_93;
    endmethod

    method ActionValue#(Struct23) cache__00__getVictim ();
        let x_1 = (victims__00);
        Struct38 x_2 = (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        (((((x_1)[(Bit#(1))'(1'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) : (Struct38 {valid :
        (Bool)'(False), data : unpack(0)})))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method Action cache__00__setVictimRq (Struct24 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(4) x_2 = ((x_0).victim_req);
        let x_3 = (victims__00);
        Struct23 x_4 =
        ((x_3)[(Bit#(1))'(1'h1)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct23 x_5 = (Struct23 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct14 {valid :
            (Bool)'(True), data : x_2}});
            victims__00 <= update (x_3, (Bit#(1))'(1'h1), x_5);
        end else begin
            Struct23 x_6 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct23 x_7 = (Struct23 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct14 {valid : (Bool)'(True), data :
                x_2}});
                victims__00 <= update (x_3, (Bit#(1))'(1'h0), x_7);
            end else begin
                Struct23 x_8 =
                ((x_3)[(Bit#(1))'(1'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct23 x_9 = (Struct23 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct14 {valid :
                    (Bool)'(True), data : x_2}});
                    victims__00 <= update (x_3, (Bit#(1))'(1'h1), x_9);
                end else begin

                end
            end
        end
    endmethod

    method ActionValue#(Bit#(4)) cache__00__releaseVictim (Bit#(64) x_0);
        let x_1 = (victims__00);
        Struct23 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victims__00 <= update (x_1, (Bit#(1))'(1'h0), unpack(0));
            Bit#(4) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct23 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victims__00 <= update (x_1, (Bit#(1))'(1'h1),
                unpack(0));
                Bit#(4) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct23 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victims__00 <= update (x_1, (Bit#(1))'(1'h0),
                    unpack(0));
                    Bit#(4) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct23 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victims__00 <= update (x_1, (Bit#(1))'(1'h1),
                        unpack(0));
                        Bit#(4) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod

    method ActionValue#(Bit#(1)) cache__00__getVictimCount ();
        let x_1 = (victims__00);
        Bit#(1) x_2 = ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((((((x_1)[(Bit#(1))'(1'h0)]).victim_valid)
        && (! ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0)))) +
        ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((Bit#(1))'(1'h0)))));
        return x_2;
    endmethod
endmodule

interface Module181;
    method Action cache__000__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct40) cache__000__infoRsValueRq ();
    method ActionValue#(Vector#(4, Bit#(64))) cache__000__valueRsLineRq
    (Struct43 x_0);
    method ActionValue#(Struct23) cache__000__getVictim ();
    method Action cache__000__setVictimRq (Struct24 x_0);
    method ActionValue#(Bit#(4)) cache__000__releaseVictim (Bit#(64) x_0);
    method ActionValue#(Bit#(1)) cache__000__getVictimCount ();
endinterface

module mkModule181#(function Action wrReq_edirRam__000__3(Struct53 _),
    function Action wrReq_edirRam__000__2(Struct53 _),
    function Action wrReq_edirRam__000__1(Struct53 _),
    function Action wrReq_edirRam__000__0(Struct53 _),
    function Action wrReq_dataRam__000(Struct52 _),
    function Action repAccess__000(Struct51 _),
    function Action wrReq_infoRam__000__7(Struct50 _),
    function Action wrReq_infoRam__000__6(Struct50 _),
    function Action wrReq_infoRam__000__5(Struct50 _),
    function Action wrReq_infoRam__000__4(Struct50 _),
    function Action wrReq_infoRam__000__3(Struct50 _),
    function Action wrReq_infoRam__000__2(Struct50 _),
    function Action wrReq_infoRam__000__1(Struct50 _),
    function Action wrReq_infoRam__000__0(Struct50 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__000(),
    function ActionValue#(Struct45) deq_cp_2__000(),
    function Action rdReq_dataRam__000(Bit#(12) _),
    function ActionValue#(Vector#(8, Bit#(8))) repGetRs__000(),
    function ActionValue#(Struct48) rdResp_edirRam__000__3(),
    function ActionValue#(Struct48) rdResp_edirRam__000__2(),
    function ActionValue#(Struct48) rdResp_edirRam__000__1(),
    function ActionValue#(Struct48) rdResp_edirRam__000__0(),
    function ActionValue#(Struct46) rdResp_infoRam__000__7(),
    function ActionValue#(Struct46) rdResp_infoRam__000__6(),
    function ActionValue#(Struct46) rdResp_infoRam__000__5(),
    function ActionValue#(Struct46) rdResp_infoRam__000__4(),
    function ActionValue#(Struct46) rdResp_infoRam__000__3(),
    function ActionValue#(Struct46) rdResp_infoRam__000__2(),
    function ActionValue#(Struct46) rdResp_infoRam__000__1(),
    function ActionValue#(Struct46) rdResp_infoRam__000__0(),
    function Action enq_cp_2__000(Struct45 _),
    function ActionValue#(Struct44) deq_cp_1__000(),
    function Action repGetRq__000(Bit#(9) _),
    function Action rdReq_edirRam__000__3(Bit#(9) _),
    function Action rdReq_edirRam__000__2(Bit#(9) _),
    function Action rdReq_edirRam__000__1(Bit#(9) _),
    function Action rdReq_edirRam__000__0(Bit#(9) _),
    function Action rdReq_infoRam__000__7(Bit#(9) _),
    function Action rdReq_infoRam__000__6(Bit#(9) _),
    function Action rdReq_infoRam__000__5(Bit#(9) _),
    function Action rdReq_infoRam__000__4(Bit#(9) _),
    function Action rdReq_infoRam__000__3(Bit#(9) _),
    function Action rdReq_infoRam__000__2(Bit#(9) _),
    function Action rdReq_infoRam__000__1(Bit#(9) _),
    function Action rdReq_infoRam__000__0(Bit#(9) _),
    function Action enq_cp_1__000(Struct44 _))
    (Module181);
    Reg#(Vector#(4, Struct23)) victims__000 <- mkReg(unpack(0));

    // No rules in this module

    method Action cache__000__infoRq (Bit#(64) x_0);
        let x_1 = (victims__000);
        Struct23 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            let x_3 <- enq_cp_1__000(Struct44 {tag : (x_0)[63:14], index :
            (x_0)[13:5], victim_found : Struct26 {valid : (Bool)'(True), data
            : (Bit#(1))'(1'h0)}});
        end else begin
            Struct23 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                let x_5 <- enq_cp_1__000(Struct44 {tag : (x_0)[63:14], index
                : (x_0)[13:5], victim_found : Struct26 {valid :
                (Bool)'(True), data : (Bit#(1))'(1'h1)}});
            end else begin
                Struct23 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    let x_7 <- enq_cp_1__000(Struct44 {tag : (x_0)[63:14],
                    index : (x_0)[13:5], victim_found : Struct26 {valid :
                    (Bool)'(True), data : (Bit#(1))'(1'h0)}});
                end else begin
                    Struct23 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        let x_9 <- enq_cp_1__000(Struct44 {tag :
                        (x_0)[63:14], index : (x_0)[13:5], victim_found :
                        Struct26 {valid : (Bool)'(True), data :
                        (Bit#(1))'(1'h1)}});
                    end else begin
                        Bit#(9) x_10 = ((x_0)[13:5]);
                        let x_11 <- rdReq_infoRam__000__0(x_10);
                        let x_12 <- rdReq_infoRam__000__1(x_10);
                        let x_13 <- rdReq_infoRam__000__2(x_10);
                        let x_14 <- rdReq_infoRam__000__3(x_10);
                        let x_15 <- rdReq_infoRam__000__4(x_10);
                        let x_16 <- rdReq_infoRam__000__5(x_10);
                        let x_17 <- rdReq_infoRam__000__6(x_10);
                        let x_18 <- rdReq_infoRam__000__7(x_10);
                        let x_19 <- rdReq_edirRam__000__0(x_10);
                        let x_20 <- rdReq_edirRam__000__1(x_10);
                        let x_21 <- rdReq_edirRam__000__2(x_10);
                        let x_22 <- rdReq_edirRam__000__3(x_10);
                        let x_23 <- repGetRq__000(x_10);
                        let x_24 <- enq_cp_1__000(Struct44 {tag :
                        (x_0)[63:14], index : (x_0)[13:5], victim_found :
                        Struct26 {valid : (Bool)'(False), data :
                        unpack(0)}});
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Struct40) cache__000__infoRsValueRq ();
        let x_1 <- deq_cp_1__000();
        Bit#(50) x_2 = ((x_1).tag);
        Bit#(9) x_3 =
        ((x_1).index);
        let x_64 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_4 = (((x_1).victim_found).data);
            let x_5 = (victims__000);
            Struct23 x_6 = ((x_5)[x_4]);
            Struct40 x_7 = (Struct40 {info_index : x_3, info_hit :
            (Bool)'(True), info_way : unpack(0), edir_hit : (Bool)'(False),
            edir_way : unpack(0), edir_slot : Struct41 {valid :
            (Bool)'(False), data : unpack(0)}, info : (x_6).victim_info});
            let x_8 <- enq_cp_2__000(Struct45 {victim_found :
            (x_1).victim_found, may_victim : unpack(0), reps :
            unpack(0)});
            x_64 = x_7;
        end else begin
            Vector#(8, Struct46) x_9 = (unpack(0));
            let x_10 <- rdResp_infoRam__000__0();
            Vector#(8, Struct46) x_11 = (update (x_9, (Bit#(3))'(3'h0),
            x_10));
            let x_12 <- rdResp_infoRam__000__1();
            Vector#(8, Struct46) x_13 = (update (x_11, (Bit#(3))'(3'h1),
            x_12));
            let x_14 <- rdResp_infoRam__000__2();
            Vector#(8, Struct46) x_15 = (update (x_13, (Bit#(3))'(3'h2),
            x_14));
            let x_16 <- rdResp_infoRam__000__3();
            Vector#(8, Struct46) x_17 = (update (x_15, (Bit#(3))'(3'h3),
            x_16));
            let x_18 <- rdResp_infoRam__000__4();
            Vector#(8, Struct46) x_19 = (update (x_17, (Bit#(3))'(3'h4),
            x_18));
            let x_20 <- rdResp_infoRam__000__5();
            Vector#(8, Struct46) x_21 = (update (x_19, (Bit#(3))'(3'h5),
            x_20));
            let x_22 <- rdResp_infoRam__000__6();
            Vector#(8, Struct46) x_23 = (update (x_21, (Bit#(3))'(3'h6),
            x_22));
            let x_24 <- rdResp_infoRam__000__7();
            Vector#(8, Struct46) x_25 = (update (x_23, (Bit#(3))'(3'h7),
            x_24));
            Struct47 x_26 = (((((x_25)[(Bit#(3))'(3'h0)]).tag) == (x_2) ?
            (Struct47 {tm_hit : (Bool)'(True), tm_way : (Bit#(3))'(3'h0),
            tm_value : ((x_25)[(Bit#(3))'(3'h0)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h1)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h1), tm_value :
            ((x_25)[(Bit#(3))'(3'h1)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h2)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h2), tm_value :
            ((x_25)[(Bit#(3))'(3'h2)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h3)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h3), tm_value :
            ((x_25)[(Bit#(3))'(3'h3)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h4)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h4), tm_value :
            ((x_25)[(Bit#(3))'(3'h4)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h5)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h5), tm_value :
            ((x_25)[(Bit#(3))'(3'h5)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h6)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h6), tm_value :
            ((x_25)[(Bit#(3))'(3'h6)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h7)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h7), tm_value :
            ((x_25)[(Bit#(3))'(3'h7)]).value}) :
            (unpack(0))))))))))))))))));
            Vector#(4, Struct48) x_27 = (unpack(0));
            let x_28 <- rdResp_edirRam__000__0();
            Vector#(4, Struct48) x_29 = (update (x_27, (Bit#(2))'(2'h0),
            x_28));
            let x_30 <- rdResp_edirRam__000__1();
            Vector#(4, Struct48) x_31 = (update (x_29, (Bit#(2))'(2'h1),
            x_30));
            let x_32 <- rdResp_edirRam__000__2();
            Vector#(4, Struct48) x_33 = (update (x_31, (Bit#(2))'(2'h2),
            x_32));
            let x_34 <- rdResp_edirRam__000__3();
            Vector#(4, Struct48) x_35 = (update (x_33, (Bit#(2))'(2'h3),
            x_34));
            Struct49 x_36 = (((((x_35)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
            (Struct49 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
            tm_value : ((x_35)[(Bit#(2))'(2'h0)]).value}) :
            (((((x_35)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct49 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
            ((x_35)[(Bit#(2))'(2'h1)]).value}) :
            (((((x_35)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct49 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
            ((x_35)[(Bit#(2))'(2'h2)]).value}) :
            (((((x_35)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct49 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
            ((x_35)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
            Struct32 x_37 = ((x_36).tm_value);
            Struct41 x_38 =
            (((((((x_35)[(Bit#(2))'(2'h0)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h0)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h0)}) :
            (((((((x_35)[(Bit#(2))'(2'h1)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h1)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h1)}) :
            (((((((x_35)[(Bit#(2))'(2'h2)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h2)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h2)}) :
            (((((((x_35)[(Bit#(2))'(2'h3)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h3)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h3)}) : (Struct41 {valid : (Bool)'(False), data :
            unpack(0)})))))))));
            let x_39 <- repGetRs__000();
            Bit#(3) x_40 = (unpack(0));
            Bit#(8) x_41 = (unpack(0));
            Bit#(3) x_42 = ((! (((x_39)[(Bit#(3))'(3'h7)]) < (x_41)) ?
            ((Bit#(3))'(3'h7)) : (x_40)));
            Bit#(8) x_43 = ((! (((x_39)[(Bit#(3))'(3'h7)]) < (x_41)) ?
            ((x_39)[(Bit#(3))'(3'h7)]) : (x_41)));
            Bit#(3) x_44 = ((! (((x_39)[(Bit#(3))'(3'h6)]) < (x_43)) ?
            ((Bit#(3))'(3'h6)) : (x_42)));
            Bit#(8) x_45 = ((! (((x_39)[(Bit#(3))'(3'h6)]) < (x_43)) ?
            ((x_39)[(Bit#(3))'(3'h6)]) : (x_43)));
            Bit#(3) x_46 = ((! (((x_39)[(Bit#(3))'(3'h5)]) < (x_45)) ?
            ((Bit#(3))'(3'h5)) : (x_44)));
            Bit#(8) x_47 = ((! (((x_39)[(Bit#(3))'(3'h5)]) < (x_45)) ?
            ((x_39)[(Bit#(3))'(3'h5)]) : (x_45)));
            Bit#(3) x_48 = ((! (((x_39)[(Bit#(3))'(3'h4)]) < (x_47)) ?
            ((Bit#(3))'(3'h4)) : (x_46)));
            Bit#(8) x_49 = ((! (((x_39)[(Bit#(3))'(3'h4)]) < (x_47)) ?
            ((x_39)[(Bit#(3))'(3'h4)]) : (x_47)));
            Bit#(3) x_50 = ((! (((x_39)[(Bit#(3))'(3'h3)]) < (x_49)) ?
            ((Bit#(3))'(3'h3)) : (x_48)));
            Bit#(8) x_51 = ((! (((x_39)[(Bit#(3))'(3'h3)]) < (x_49)) ?
            ((x_39)[(Bit#(3))'(3'h3)]) : (x_49)));
            Bit#(3) x_52 = ((! (((x_39)[(Bit#(3))'(3'h2)]) < (x_51)) ?
            ((Bit#(3))'(3'h2)) : (x_50)));
            Bit#(8) x_53 = ((! (((x_39)[(Bit#(3))'(3'h2)]) < (x_51)) ?
            ((x_39)[(Bit#(3))'(3'h2)]) : (x_51)));
            Bit#(3) x_54 = ((! (((x_39)[(Bit#(3))'(3'h1)]) < (x_53)) ?
            ((Bit#(3))'(3'h1)) : (x_52)));
            Bit#(8) x_55 = ((! (((x_39)[(Bit#(3))'(3'h1)]) < (x_53)) ?
            ((x_39)[(Bit#(3))'(3'h1)]) : (x_53)));
            Bit#(3) x_56 = ((! (((x_39)[(Bit#(3))'(3'h0)]) < (x_55)) ?
            ((Bit#(3))'(3'h0)) : (x_54)));
            Bit#(8) x_57 = ((! (((x_39)[(Bit#(3))'(3'h0)]) < (x_55)) ?
            ((x_39)[(Bit#(3))'(3'h0)]) : (x_55)));
            Struct40 x_58 = (Struct40 {info_index : x_3, info_hit :
            (x_26).tm_hit, info_way : (x_26).tm_way, edir_hit :
            (x_36).tm_hit, edir_way : (x_36).tm_way, edir_slot : x_38, info :
            ((x_26).tm_hit ? ((x_26).tm_value) : (Struct11 {mesi_owned :
            (Bool)'(False), mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
            (x_37).mesi_edir_st, mesi_dir_sharers :
            (x_37).mesi_edir_sharers}))});
            Struct46 x_59 = ((x_25)[x_56]);
            Bit#(50) x_60 = ((x_59).tag);
            Struct11 x_61 = ((x_59).value);
            let x_62 <- enq_cp_2__000(Struct45 {victim_found : Struct26
            {valid : (Bool)'(False), data : unpack(0)}, may_victim : Struct28
            {mv_addr : {(x_60),({(x_3),((Bit#(5))'(5'h0))})}, mv_info :
            x_61}, reps : x_39});
            let x_63 <- rdReq_dataRam__000({(((x_26).tm_hit ? ((x_26).tm_way)
            : (x_56))),(x_3)});
            x_64 = x_58;
        end
        return x_64;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__000__valueRsLineRq
    (Struct43 x_0);
        let x_1 <- deq_cp_2__000();
        let x_2 =
        (victims__000);
        let x_61 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_3 = (((x_1).victim_found).data);
            Struct23 x_4 = ((x_2)[x_3]);
            Struct23 x_5 = (Struct23 {victim_valid : (Bool)'(True),
            victim_addr : (x_4).victim_addr, victim_info : ((x_0).info_write
            ? ((x_0).info) : ((x_4).victim_info)), victim_value :
            ((x_0).value_write ? ((x_0).value) : ((x_4).victim_value)),
            victim_req : (x_4).victim_req});
            victims__000 <= update (x_2, x_3, x_5);
            x_61 = (x_4).victim_value;
        end else begin
            let x_6 <- rdResp_dataRam__000();
            Bit#(64) x_7 = ((x_0).addr);
            Bit#(9) x_8 = ((x_7)[13:5]);
            Bit#(3) x_9 = ((x_0).info_way);
            Struct11 x_10 = ((x_0).info);
            Bool x_11 = ((! ((x_10).mesi_owned)) && (((x_10).mesi_status) ==
            ((Bit#(3))'(3'h1))));
            if ((((x_0).info_hit) || (! (x_11))) || ((! ((x_0).edir_hit)) &&
                (x_11)))
                begin
                if ((x_0).info_write) begin
                    Struct50 x_12 = (Struct50 {addr : x_8, datain : Struct46
                    {tag : (x_7)[63:14], value :
                    x_10}});
                    if ((x_9) == ((Bit#(3))'(3'h0))) begin
                        let x_13 <- wrReq_infoRam__000__0(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h1))) begin
                        let x_15 <- wrReq_infoRam__000__1(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h2))) begin
                        let x_17 <- wrReq_infoRam__000__2(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h3))) begin
                        let x_19 <- wrReq_infoRam__000__3(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h4))) begin
                        let x_21 <- wrReq_infoRam__000__4(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h5))) begin
                        let x_23 <- wrReq_infoRam__000__5(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h6))) begin
                        let x_25 <- wrReq_infoRam__000__6(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h7))) begin
                        let x_27 <- wrReq_infoRam__000__7(x_12);
                    end else begin

                    end
                    Struct28 x_29 = ((x_1).may_victim);
                    Struct26 x_30 = ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid
                    ? ((((x_2)[(Bit#(1))'(1'h0)]).victim_valid ?
                    ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid ? (Struct26
                    {valid : (Bool)'(False), data : unpack(0)}) : (Struct26
                    {valid : (Bool)'(True), data : (Bit#(1))'(1'h1)}))) :
                    (Struct26 {valid : (Bool)'(True), data :
                    (Bit#(1))'(1'h0)}))) : (Struct26 {valid : (Bool)'(True),
                    data : (Bit#(1))'(1'h1)})));
                    Bit#(1) x_31 = ((x_30).data);
                    victims__000 <= update (x_2, x_31, Struct23 {victim_valid
                    : (Bool)'(True), victim_addr : (x_29).mv_addr,
                    victim_info : (x_29).mv_info, victim_value : x_6,
                    victim_req : Struct14 {valid : (Bool)'(False), data :
                    unpack(0)}});
                    let x_32 <- repAccess__000(Struct51 {acc_type :
                    ((((x_10).mesi_dir_st) == ((Bit#(3))'(3'h0))) ||
                    (((x_10).mesi_dir_st) == ((Bit#(3))'(3'h1))) ?
                    ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))), acc_reps :
                    (x_1).reps, acc_index : x_8, acc_way : x_9});
                end else begin

                end
                if ((x_0).value_write) begin
                    Struct52 x_34 = (Struct52 {addr : {(x_9),((x_7)[13:5])},
                    datain : (x_0).value});
                    let x_35 <- wrReq_dataRam__000(x_34);
                end else begin

                end
            end else begin

            end
            if (((x_0).info_write) && ((x_0).edir_hit)) begin
                Bit#(2) x_38 = ((x_0).edir_way);
                Struct53 x_39 = (Struct53 {addr : (x_7)[13:5], datain :
                Struct48 {tag : (x_7)[63:14], value : (x_11 ? (Struct32
                {mesi_edir_st : (x_10).mesi_dir_st, mesi_edir_sharers :
                (x_10).mesi_dir_sharers}) :
                (unpack(0)))}});
                if ((x_38) == ((Bit#(2))'(2'h0))) begin
                    let x_40 <- wrReq_edirRam__000__0(x_39);
                end else begin

                end
                if ((x_38) == ((Bit#(2))'(2'h1))) begin
                    let x_42 <- wrReq_edirRam__000__1(x_39);
                end else begin

                end
                if ((x_38) == ((Bit#(2))'(2'h2))) begin
                    let x_44 <- wrReq_edirRam__000__2(x_39);
                end else begin

                end
                if ((x_38) == ((Bit#(2))'(2'h3))) begin
                    let x_46 <- wrReq_edirRam__000__3(x_39);
                end else begin

                end
            end else begin
                Struct41 x_48 =
                ((x_0).edir_slot);
                if (((! ((x_0).edir_hit)) && ((x_48).valid)) && (x_11))
                    begin
                    Bit#(2) x_49 = ((x_48).data);
                    Struct53 x_50 = (Struct53 {addr : (x_7)[13:5], datain :
                    Struct48 {tag : (x_7)[63:14], value : Struct32
                    {mesi_edir_st : (x_10).mesi_dir_st, mesi_edir_sharers :
                    (x_10).mesi_dir_sharers}}});
                    if ((x_49) == ((Bit#(2))'(2'h0))) begin
                        let x_51 <- wrReq_edirRam__000__0(x_50);
                    end else begin

                    end
                    if ((x_49) == ((Bit#(2))'(2'h1))) begin
                        let x_53 <- wrReq_edirRam__000__1(x_50);
                    end else begin

                    end
                    if ((x_49) == ((Bit#(2))'(2'h2))) begin
                        let x_55 <- wrReq_edirRam__000__2(x_50);
                    end else begin

                    end
                    if ((x_49) == ((Bit#(2))'(2'h3))) begin
                        let x_57 <- wrReq_edirRam__000__3(x_50);
                    end else begin

                    end
                end else begin

                end
            end
            x_61 = x_6;
        end
        return x_61;
    endmethod

    method ActionValue#(Struct23) cache__000__getVictim ();
        let x_1 = (victims__000);
        Struct38 x_2 = (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        (((((x_1)[(Bit#(1))'(1'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) : (Struct38 {valid :
        (Bool)'(False), data : unpack(0)})))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method Action cache__000__setVictimRq (Struct24 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(4) x_2 = ((x_0).victim_req);
        let x_3 = (victims__000);
        Struct23 x_4 =
        ((x_3)[(Bit#(1))'(1'h1)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct23 x_5 = (Struct23 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct14 {valid :
            (Bool)'(True), data : x_2}});
            victims__000 <= update (x_3, (Bit#(1))'(1'h1), x_5);
        end else begin
            Struct23 x_6 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct23 x_7 = (Struct23 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct14 {valid : (Bool)'(True), data :
                x_2}});
                victims__000 <= update (x_3, (Bit#(1))'(1'h0), x_7);
            end else begin
                Struct23 x_8 =
                ((x_3)[(Bit#(1))'(1'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct23 x_9 = (Struct23 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct14 {valid :
                    (Bool)'(True), data : x_2}});
                    victims__000 <= update (x_3, (Bit#(1))'(1'h1), x_9);
                end else begin

                end
            end
        end
    endmethod

    method ActionValue#(Bit#(4)) cache__000__releaseVictim (Bit#(64) x_0);
        let x_1 = (victims__000);
        Struct23 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victims__000 <= update (x_1, (Bit#(1))'(1'h0), unpack(0));
            Bit#(4) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct23 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victims__000 <= update (x_1, (Bit#(1))'(1'h1),
                unpack(0));
                Bit#(4) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct23 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victims__000 <= update (x_1, (Bit#(1))'(1'h0),
                    unpack(0));
                    Bit#(4) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct23 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victims__000 <= update (x_1, (Bit#(1))'(1'h1),
                        unpack(0));
                        Bit#(4) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod

    method ActionValue#(Bit#(1)) cache__000__getVictimCount ();
        let x_1 = (victims__000);
        Bit#(1) x_2 = ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((((((x_1)[(Bit#(1))'(1'h0)]).victim_valid)
        && (! ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0)))) +
        ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((Bit#(1))'(1'h0)))));
        return x_2;
    endmethod
endmodule

interface Module182;
    method Action cache__0000__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct60) cache__0000__infoRsValueRq ();
    method ActionValue#(Vector#(4, Bit#(64))) cache__0000__valueRsLineRq
    (Struct64 x_0);
    method ActionValue#(Struct66) cache__0000__getVictim ();
    method Action cache__0000__setVictimRq (Struct67 x_0);
    method ActionValue#(Bit#(3)) cache__0000__releaseVictim (Bit#(64) x_0);
    method ActionValue#(Bit#(1)) cache__0000__getVictimCount ();
endinterface

module mkModule182#(function Action repAccess__0000(Struct74 _),
    function Action wrReq_dataRam__0000(Struct73 _),
    function Action wrReq_infoRam__0000__3(Struct72 _),
    function Action wrReq_infoRam__0000__2(Struct72 _),
    function Action wrReq_infoRam__0000__1(Struct72 _),
    function Action wrReq_infoRam__0000__0(Struct72 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0000(),
    function ActionValue#(Struct69) deq_cp_2__0000(),
    function Action rdReq_dataRam__0000(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__0000(),
    function ActionValue#(Struct70) rdResp_infoRam__0000__3(),
    function ActionValue#(Struct70) rdResp_infoRam__0000__2(),
    function ActionValue#(Struct70) rdResp_infoRam__0000__1(),
    function ActionValue#(Struct70) rdResp_infoRam__0000__0(),
    function Action enq_cp_2__0000(Struct69 _),
    function ActionValue#(Struct68) deq_cp_1__0000(),
    function Action repGetRq__0000(Bit#(8) _),
    function Action rdReq_infoRam__0000__3(Bit#(8) _),
    function Action rdReq_infoRam__0000__2(Bit#(8) _),
    function Action rdReq_infoRam__0000__1(Bit#(8) _),
    function Action rdReq_infoRam__0000__0(Bit#(8) _),
    function Action enq_cp_1__0000(Struct68 _))
    (Module182);
    Reg#(Vector#(4, Struct66)) victims__0000 <- mkReg(unpack(0));

    // No rules in this module

    method Action cache__0000__infoRq (Bit#(64) x_0);
        let x_1 = (victims__0000);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            let x_3 <- enq_cp_1__0000(Struct68 {tag : (x_0)[63:13], index :
            (x_0)[12:5], victim_found : Struct26 {valid : (Bool)'(True), data
            : (Bit#(1))'(1'h0)}});
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                let x_5 <- enq_cp_1__0000(Struct68 {tag : (x_0)[63:13], index
                : (x_0)[12:5], victim_found : Struct26 {valid :
                (Bool)'(True), data : (Bit#(1))'(1'h1)}});
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    let x_7 <- enq_cp_1__0000(Struct68 {tag : (x_0)[63:13],
                    index : (x_0)[12:5], victim_found : Struct26 {valid :
                    (Bool)'(True), data : (Bit#(1))'(1'h0)}});
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        let x_9 <- enq_cp_1__0000(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(True), data :
                        (Bit#(1))'(1'h1)}});
                    end else begin
                        Bit#(8) x_10 = ((x_0)[12:5]);
                        let x_11 <- rdReq_infoRam__0000__0(x_10);
                        let x_12 <- rdReq_infoRam__0000__1(x_10);
                        let x_13 <- rdReq_infoRam__0000__2(x_10);
                        let x_14 <- rdReq_infoRam__0000__3(x_10);
                        let x_15 <- repGetRq__0000(x_10);
                        let x_16 <- enq_cp_1__0000(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(False), data :
                        unpack(0)}});
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Struct60) cache__0000__infoRsValueRq ();
        let x_1 <- deq_cp_1__0000();
        Bit#(51) x_2 = ((x_1).tag);
        Bit#(8) x_3 =
        ((x_1).index);
        let x_36 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_4 = (((x_1).victim_found).data);
            let x_5 = (victims__0000);
            Struct66 x_6 = ((x_5)[x_4]);
            Struct60 x_7 = (Struct60 {info_index : x_3, info_hit :
            (Bool)'(True), info_way : unpack(0), edir_hit : (Bool)'(False),
            edir_way : unpack(0), edir_slot : Struct61 {valid :
            (Bool)'(False), data : unpack(0)}, info : (x_6).victim_info});
            let x_8 <- enq_cp_2__0000(Struct69 {victim_found :
            (x_1).victim_found, may_victim : unpack(0), reps :
            unpack(0)});
            x_36 = x_7;
        end else begin
            Vector#(4, Struct70) x_9 = (unpack(0));
            let x_10 <- rdResp_infoRam__0000__0();
            Vector#(4, Struct70) x_11 = (update (x_9, (Bit#(2))'(2'h0),
            x_10));
            let x_12 <- rdResp_infoRam__0000__1();
            Vector#(4, Struct70) x_13 = (update (x_11, (Bit#(2))'(2'h1),
            x_12));
            let x_14 <- rdResp_infoRam__0000__2();
            Vector#(4, Struct70) x_15 = (update (x_13, (Bit#(2))'(2'h2),
            x_14));
            let x_16 <- rdResp_infoRam__0000__3();
            Vector#(4, Struct70) x_17 = (update (x_15, (Bit#(2))'(2'h3),
            x_16));
            Struct71 x_18 = (((((x_17)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
            (Struct71 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
            tm_value : ((x_17)[(Bit#(2))'(2'h0)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
            ((x_17)[(Bit#(2))'(2'h1)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
            ((x_17)[(Bit#(2))'(2'h2)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
            ((x_17)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
            let x_19 <- repGetRs__0000();
            Bit#(2) x_20 = (unpack(0));
            Bit#(8) x_21 = (unpack(0));
            Bit#(2) x_22 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((Bit#(2))'(2'h3)) : (x_20)));
            Bit#(8) x_23 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((x_19)[(Bit#(2))'(2'h3)]) : (x_21)));
            Bit#(2) x_24 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((Bit#(2))'(2'h2)) : (x_22)));
            Bit#(8) x_25 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((x_19)[(Bit#(2))'(2'h2)]) : (x_23)));
            Bit#(2) x_26 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((Bit#(2))'(2'h1)) : (x_24)));
            Bit#(8) x_27 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((x_19)[(Bit#(2))'(2'h1)]) : (x_25)));
            Bit#(2) x_28 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((Bit#(2))'(2'h0)) : (x_26)));
            Bit#(8) x_29 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((x_19)[(Bit#(2))'(2'h0)]) : (x_27)));
            Struct60 x_30 = (Struct60 {info_index : x_3, info_hit :
            (x_18).tm_hit, info_way : (x_18).tm_way, edir_hit : unpack(0),
            edir_way : unpack(0), edir_slot : unpack(0), info :
            (x_18).tm_value});
            Struct70 x_31 = ((x_17)[x_28]);
            Bit#(51) x_32 = ((x_31).tag);
            Struct11 x_33 = ((x_31).value);
            let x_34 <- enq_cp_2__0000(Struct69 {victim_found : Struct26
            {valid : (Bool)'(False), data : unpack(0)}, may_victim : Struct28
            {mv_addr : {(x_32),({(x_3),((Bit#(5))'(5'h0))})}, mv_info :
            x_33}, reps : x_19});
            let x_35 <- rdReq_dataRam__0000({(((x_18).tm_hit ?
            ((x_18).tm_way) : (x_28))),(x_3)});
            x_36 = x_30;
        end
        return x_36;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__0000__valueRsLineRq
    (Struct64 x_0);
        let x_1 <- deq_cp_2__0000();
        let x_2 =
        (victims__0000);
        let x_29 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_3 = (((x_1).victim_found).data);
            Struct66 x_4 = ((x_2)[x_3]);
            Struct66 x_5 = (Struct66 {victim_valid : (Bool)'(True),
            victim_addr : (x_4).victim_addr, victim_info : ((x_0).info_write
            ? ((x_0).info) : ((x_4).victim_info)), victim_value :
            ((x_0).value_write ? ((x_0).value) : ((x_4).victim_value)),
            victim_req : (x_4).victim_req});
            victims__0000 <= update (x_2, x_3, x_5);
            x_29 = (x_4).victim_value;
        end else begin
            let x_6 <- rdResp_dataRam__0000();
            Bit#(64) x_7 = ((x_0).addr);
            Bit#(8) x_8 = ((x_7)[12:5]);
            Bit#(2) x_9 = ((x_0).info_way);
            Struct11 x_10 =
            ((x_0).info);
            if ((x_0).info_write) begin
                Struct72 x_11 = (Struct72 {addr : x_8, datain : Struct70 {tag
                : (x_7)[63:13], value :
                x_10}});
                if ((x_9) == ((Bit#(2))'(2'h0))) begin
                    let x_12 <- wrReq_infoRam__0000__0(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h1))) begin
                    let x_14 <- wrReq_infoRam__0000__1(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h2))) begin
                    let x_16 <- wrReq_infoRam__0000__2(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h3))) begin
                    let x_18 <- wrReq_infoRam__0000__3(x_11);
                end else begin

                end
                if ((x_0).value_write) begin
                    Struct73 x_20 = (Struct73 {addr : {(x_9),((x_7)[12:5])},
                    datain : (x_0).value});
                    let x_21 <- wrReq_dataRam__0000(x_20);
                end else begin

                end
                if (! ((x_0).info_hit)) begin
                    Struct28 x_23 = ((x_1).may_victim);
                    Struct26 x_24 = ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid
                    ? ((((x_2)[(Bit#(1))'(1'h0)]).victim_valid ?
                    ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid ? (Struct26
                    {valid : (Bool)'(False), data : unpack(0)}) : (Struct26
                    {valid : (Bool)'(True), data : (Bit#(1))'(1'h1)}))) :
                    (Struct26 {valid : (Bool)'(True), data :
                    (Bit#(1))'(1'h0)}))) : (Struct26 {valid : (Bool)'(True),
                    data : (Bit#(1))'(1'h1)})));
                    Bit#(1) x_25 = ((x_24).data);
                    victims__0000 <= update (x_2, x_25, Struct66
                    {victim_valid : (Bool)'(True), victim_addr :
                    (x_23).mv_addr, victim_info : (x_23).mv_info,
                    victim_value : x_6, victim_req : Struct10 {valid :
                    (Bool)'(False), data : unpack(0)}});
                end else begin

                end
                let x_27 <- repAccess__0000(Struct74 {acc_type :
                ((((x_10).mesi_dir_st) == ((Bit#(3))'(3'h0))) ||
                (((x_10).mesi_dir_st) == ((Bit#(3))'(3'h1))) ?
                ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))), acc_reps :
                (x_1).reps, acc_index : x_8, acc_way : x_9});
            end else begin

            end
            x_29 = x_6;
        end
        return x_29;
    endmethod

    method ActionValue#(Struct66) cache__0000__getVictim ();
        let x_1 = (victims__0000);
        Struct75 x_2 = (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        (((((x_1)[(Bit#(1))'(1'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) : (Struct75 {valid :
        (Bool)'(False), data : unpack(0)})))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method Action cache__0000__setVictimRq (Struct67 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victims__0000);
        Struct66 x_4 =
        ((x_3)[(Bit#(1))'(1'h1)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct66 x_5 = (Struct66 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct10 {valid :
            (Bool)'(True), data : x_2}});
            victims__0000 <= update (x_3, (Bit#(1))'(1'h1), x_5);
        end else begin
            Struct66 x_6 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct66 x_7 = (Struct66 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct10 {valid : (Bool)'(True), data :
                x_2}});
                victims__0000 <= update (x_3, (Bit#(1))'(1'h0), x_7);
            end else begin
                Struct66 x_8 =
                ((x_3)[(Bit#(1))'(1'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct66 x_9 = (Struct66 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct10 {valid :
                    (Bool)'(True), data : x_2}});
                    victims__0000 <= update (x_3, (Bit#(1))'(1'h1), x_9);
                end else begin

                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) cache__0000__releaseVictim (Bit#(64) x_0);
        let x_1 = (victims__0000);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victims__0000 <= update (x_1, (Bit#(1))'(1'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victims__0000 <= update (x_1, (Bit#(1))'(1'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victims__0000 <= update (x_1, (Bit#(1))'(1'h0),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victims__0000 <= update (x_1, (Bit#(1))'(1'h1),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod

    method ActionValue#(Bit#(1)) cache__0000__getVictimCount ();
        let x_1 = (victims__0000);
        Bit#(1) x_2 = ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((((((x_1)[(Bit#(1))'(1'h0)]).victim_valid)
        && (! ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0)))) +
        ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((Bit#(1))'(1'h0)))));
        return x_2;
    endmethod
endmodule

interface Module183;
    method Action cache__0001__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct60) cache__0001__infoRsValueRq ();
    method ActionValue#(Vector#(4, Bit#(64))) cache__0001__valueRsLineRq
    (Struct64 x_0);
    method ActionValue#(Struct66) cache__0001__getVictim ();
    method Action cache__0001__setVictimRq (Struct67 x_0);
    method ActionValue#(Bit#(3)) cache__0001__releaseVictim (Bit#(64) x_0);
    method ActionValue#(Bit#(1)) cache__0001__getVictimCount ();
endinterface

module mkModule183#(function Action repAccess__0001(Struct74 _),
    function Action wrReq_dataRam__0001(Struct73 _),
    function Action wrReq_infoRam__0001__3(Struct72 _),
    function Action wrReq_infoRam__0001__2(Struct72 _),
    function Action wrReq_infoRam__0001__1(Struct72 _),
    function Action wrReq_infoRam__0001__0(Struct72 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0001(),
    function ActionValue#(Struct69) deq_cp_2__0001(),
    function Action rdReq_dataRam__0001(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__0001(),
    function ActionValue#(Struct70) rdResp_infoRam__0001__3(),
    function ActionValue#(Struct70) rdResp_infoRam__0001__2(),
    function ActionValue#(Struct70) rdResp_infoRam__0001__1(),
    function ActionValue#(Struct70) rdResp_infoRam__0001__0(),
    function Action enq_cp_2__0001(Struct69 _),
    function ActionValue#(Struct68) deq_cp_1__0001(),
    function Action repGetRq__0001(Bit#(8) _),
    function Action rdReq_infoRam__0001__3(Bit#(8) _),
    function Action rdReq_infoRam__0001__2(Bit#(8) _),
    function Action rdReq_infoRam__0001__1(Bit#(8) _),
    function Action rdReq_infoRam__0001__0(Bit#(8) _),
    function Action enq_cp_1__0001(Struct68 _))
    (Module183);
    Reg#(Vector#(4, Struct66)) victims__0001 <- mkReg(unpack(0));

    // No rules in this module

    method Action cache__0001__infoRq (Bit#(64) x_0);
        let x_1 = (victims__0001);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            let x_3 <- enq_cp_1__0001(Struct68 {tag : (x_0)[63:13], index :
            (x_0)[12:5], victim_found : Struct26 {valid : (Bool)'(True), data
            : (Bit#(1))'(1'h0)}});
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                let x_5 <- enq_cp_1__0001(Struct68 {tag : (x_0)[63:13], index
                : (x_0)[12:5], victim_found : Struct26 {valid :
                (Bool)'(True), data : (Bit#(1))'(1'h1)}});
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    let x_7 <- enq_cp_1__0001(Struct68 {tag : (x_0)[63:13],
                    index : (x_0)[12:5], victim_found : Struct26 {valid :
                    (Bool)'(True), data : (Bit#(1))'(1'h0)}});
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        let x_9 <- enq_cp_1__0001(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(True), data :
                        (Bit#(1))'(1'h1)}});
                    end else begin
                        Bit#(8) x_10 = ((x_0)[12:5]);
                        let x_11 <- rdReq_infoRam__0001__0(x_10);
                        let x_12 <- rdReq_infoRam__0001__1(x_10);
                        let x_13 <- rdReq_infoRam__0001__2(x_10);
                        let x_14 <- rdReq_infoRam__0001__3(x_10);
                        let x_15 <- repGetRq__0001(x_10);
                        let x_16 <- enq_cp_1__0001(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(False), data :
                        unpack(0)}});
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Struct60) cache__0001__infoRsValueRq ();
        let x_1 <- deq_cp_1__0001();
        Bit#(51) x_2 = ((x_1).tag);
        Bit#(8) x_3 =
        ((x_1).index);
        let x_36 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_4 = (((x_1).victim_found).data);
            let x_5 = (victims__0001);
            Struct66 x_6 = ((x_5)[x_4]);
            Struct60 x_7 = (Struct60 {info_index : x_3, info_hit :
            (Bool)'(True), info_way : unpack(0), edir_hit : (Bool)'(False),
            edir_way : unpack(0), edir_slot : Struct61 {valid :
            (Bool)'(False), data : unpack(0)}, info : (x_6).victim_info});
            let x_8 <- enq_cp_2__0001(Struct69 {victim_found :
            (x_1).victim_found, may_victim : unpack(0), reps :
            unpack(0)});
            x_36 = x_7;
        end else begin
            Vector#(4, Struct70) x_9 = (unpack(0));
            let x_10 <- rdResp_infoRam__0001__0();
            Vector#(4, Struct70) x_11 = (update (x_9, (Bit#(2))'(2'h0),
            x_10));
            let x_12 <- rdResp_infoRam__0001__1();
            Vector#(4, Struct70) x_13 = (update (x_11, (Bit#(2))'(2'h1),
            x_12));
            let x_14 <- rdResp_infoRam__0001__2();
            Vector#(4, Struct70) x_15 = (update (x_13, (Bit#(2))'(2'h2),
            x_14));
            let x_16 <- rdResp_infoRam__0001__3();
            Vector#(4, Struct70) x_17 = (update (x_15, (Bit#(2))'(2'h3),
            x_16));
            Struct71 x_18 = (((((x_17)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
            (Struct71 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
            tm_value : ((x_17)[(Bit#(2))'(2'h0)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
            ((x_17)[(Bit#(2))'(2'h1)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
            ((x_17)[(Bit#(2))'(2'h2)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
            ((x_17)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
            let x_19 <- repGetRs__0001();
            Bit#(2) x_20 = (unpack(0));
            Bit#(8) x_21 = (unpack(0));
            Bit#(2) x_22 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((Bit#(2))'(2'h3)) : (x_20)));
            Bit#(8) x_23 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((x_19)[(Bit#(2))'(2'h3)]) : (x_21)));
            Bit#(2) x_24 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((Bit#(2))'(2'h2)) : (x_22)));
            Bit#(8) x_25 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((x_19)[(Bit#(2))'(2'h2)]) : (x_23)));
            Bit#(2) x_26 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((Bit#(2))'(2'h1)) : (x_24)));
            Bit#(8) x_27 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((x_19)[(Bit#(2))'(2'h1)]) : (x_25)));
            Bit#(2) x_28 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((Bit#(2))'(2'h0)) : (x_26)));
            Bit#(8) x_29 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((x_19)[(Bit#(2))'(2'h0)]) : (x_27)));
            Struct60 x_30 = (Struct60 {info_index : x_3, info_hit :
            (x_18).tm_hit, info_way : (x_18).tm_way, edir_hit : unpack(0),
            edir_way : unpack(0), edir_slot : unpack(0), info :
            (x_18).tm_value});
            Struct70 x_31 = ((x_17)[x_28]);
            Bit#(51) x_32 = ((x_31).tag);
            Struct11 x_33 = ((x_31).value);
            let x_34 <- enq_cp_2__0001(Struct69 {victim_found : Struct26
            {valid : (Bool)'(False), data : unpack(0)}, may_victim : Struct28
            {mv_addr : {(x_32),({(x_3),((Bit#(5))'(5'h0))})}, mv_info :
            x_33}, reps : x_19});
            let x_35 <- rdReq_dataRam__0001({(((x_18).tm_hit ?
            ((x_18).tm_way) : (x_28))),(x_3)});
            x_36 = x_30;
        end
        return x_36;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__0001__valueRsLineRq
    (Struct64 x_0);
        let x_1 <- deq_cp_2__0001();
        let x_2 =
        (victims__0001);
        let x_29 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_3 = (((x_1).victim_found).data);
            Struct66 x_4 = ((x_2)[x_3]);
            Struct66 x_5 = (Struct66 {victim_valid : (Bool)'(True),
            victim_addr : (x_4).victim_addr, victim_info : ((x_0).info_write
            ? ((x_0).info) : ((x_4).victim_info)), victim_value :
            ((x_0).value_write ? ((x_0).value) : ((x_4).victim_value)),
            victim_req : (x_4).victim_req});
            victims__0001 <= update (x_2, x_3, x_5);
            x_29 = (x_4).victim_value;
        end else begin
            let x_6 <- rdResp_dataRam__0001();
            Bit#(64) x_7 = ((x_0).addr);
            Bit#(8) x_8 = ((x_7)[12:5]);
            Bit#(2) x_9 = ((x_0).info_way);
            Struct11 x_10 =
            ((x_0).info);
            if ((x_0).info_write) begin
                Struct72 x_11 = (Struct72 {addr : x_8, datain : Struct70 {tag
                : (x_7)[63:13], value :
                x_10}});
                if ((x_9) == ((Bit#(2))'(2'h0))) begin
                    let x_12 <- wrReq_infoRam__0001__0(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h1))) begin
                    let x_14 <- wrReq_infoRam__0001__1(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h2))) begin
                    let x_16 <- wrReq_infoRam__0001__2(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h3))) begin
                    let x_18 <- wrReq_infoRam__0001__3(x_11);
                end else begin

                end
                if ((x_0).value_write) begin
                    Struct73 x_20 = (Struct73 {addr : {(x_9),((x_7)[12:5])},
                    datain : (x_0).value});
                    let x_21 <- wrReq_dataRam__0001(x_20);
                end else begin

                end
                if (! ((x_0).info_hit)) begin
                    Struct28 x_23 = ((x_1).may_victim);
                    Struct26 x_24 = ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid
                    ? ((((x_2)[(Bit#(1))'(1'h0)]).victim_valid ?
                    ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid ? (Struct26
                    {valid : (Bool)'(False), data : unpack(0)}) : (Struct26
                    {valid : (Bool)'(True), data : (Bit#(1))'(1'h1)}))) :
                    (Struct26 {valid : (Bool)'(True), data :
                    (Bit#(1))'(1'h0)}))) : (Struct26 {valid : (Bool)'(True),
                    data : (Bit#(1))'(1'h1)})));
                    Bit#(1) x_25 = ((x_24).data);
                    victims__0001 <= update (x_2, x_25, Struct66
                    {victim_valid : (Bool)'(True), victim_addr :
                    (x_23).mv_addr, victim_info : (x_23).mv_info,
                    victim_value : x_6, victim_req : Struct10 {valid :
                    (Bool)'(False), data : unpack(0)}});
                end else begin

                end
                let x_27 <- repAccess__0001(Struct74 {acc_type :
                ((((x_10).mesi_dir_st) == ((Bit#(3))'(3'h0))) ||
                (((x_10).mesi_dir_st) == ((Bit#(3))'(3'h1))) ?
                ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))), acc_reps :
                (x_1).reps, acc_index : x_8, acc_way : x_9});
            end else begin

            end
            x_29 = x_6;
        end
        return x_29;
    endmethod

    method ActionValue#(Struct66) cache__0001__getVictim ();
        let x_1 = (victims__0001);
        Struct75 x_2 = (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        (((((x_1)[(Bit#(1))'(1'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) : (Struct75 {valid :
        (Bool)'(False), data : unpack(0)})))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method Action cache__0001__setVictimRq (Struct67 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victims__0001);
        Struct66 x_4 =
        ((x_3)[(Bit#(1))'(1'h1)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct66 x_5 = (Struct66 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct10 {valid :
            (Bool)'(True), data : x_2}});
            victims__0001 <= update (x_3, (Bit#(1))'(1'h1), x_5);
        end else begin
            Struct66 x_6 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct66 x_7 = (Struct66 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct10 {valid : (Bool)'(True), data :
                x_2}});
                victims__0001 <= update (x_3, (Bit#(1))'(1'h0), x_7);
            end else begin
                Struct66 x_8 =
                ((x_3)[(Bit#(1))'(1'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct66 x_9 = (Struct66 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct10 {valid :
                    (Bool)'(True), data : x_2}});
                    victims__0001 <= update (x_3, (Bit#(1))'(1'h1), x_9);
                end else begin

                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) cache__0001__releaseVictim (Bit#(64) x_0);
        let x_1 = (victims__0001);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victims__0001 <= update (x_1, (Bit#(1))'(1'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victims__0001 <= update (x_1, (Bit#(1))'(1'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victims__0001 <= update (x_1, (Bit#(1))'(1'h0),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victims__0001 <= update (x_1, (Bit#(1))'(1'h1),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod

    method ActionValue#(Bit#(1)) cache__0001__getVictimCount ();
        let x_1 = (victims__0001);
        Bit#(1) x_2 = ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((((((x_1)[(Bit#(1))'(1'h0)]).victim_valid)
        && (! ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0)))) +
        ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((Bit#(1))'(1'h0)))));
        return x_2;
    endmethod
endmodule

interface Module184;
    method Action cache__001__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct40) cache__001__infoRsValueRq ();
    method ActionValue#(Vector#(4, Bit#(64))) cache__001__valueRsLineRq
    (Struct43 x_0);
    method ActionValue#(Struct23) cache__001__getVictim ();
    method Action cache__001__setVictimRq (Struct24 x_0);
    method ActionValue#(Bit#(4)) cache__001__releaseVictim (Bit#(64) x_0);
    method ActionValue#(Bit#(1)) cache__001__getVictimCount ();
endinterface

module mkModule184#(function Action wrReq_edirRam__001__3(Struct53 _),
    function Action wrReq_edirRam__001__2(Struct53 _),
    function Action wrReq_edirRam__001__1(Struct53 _),
    function Action wrReq_edirRam__001__0(Struct53 _),
    function Action wrReq_dataRam__001(Struct52 _),
    function Action repAccess__001(Struct51 _),
    function Action wrReq_infoRam__001__7(Struct50 _),
    function Action wrReq_infoRam__001__6(Struct50 _),
    function Action wrReq_infoRam__001__5(Struct50 _),
    function Action wrReq_infoRam__001__4(Struct50 _),
    function Action wrReq_infoRam__001__3(Struct50 _),
    function Action wrReq_infoRam__001__2(Struct50 _),
    function Action wrReq_infoRam__001__1(Struct50 _),
    function Action wrReq_infoRam__001__0(Struct50 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__001(),
    function ActionValue#(Struct45) deq_cp_2__001(),
    function Action rdReq_dataRam__001(Bit#(12) _),
    function ActionValue#(Vector#(8, Bit#(8))) repGetRs__001(),
    function ActionValue#(Struct48) rdResp_edirRam__001__3(),
    function ActionValue#(Struct48) rdResp_edirRam__001__2(),
    function ActionValue#(Struct48) rdResp_edirRam__001__1(),
    function ActionValue#(Struct48) rdResp_edirRam__001__0(),
    function ActionValue#(Struct46) rdResp_infoRam__001__7(),
    function ActionValue#(Struct46) rdResp_infoRam__001__6(),
    function ActionValue#(Struct46) rdResp_infoRam__001__5(),
    function ActionValue#(Struct46) rdResp_infoRam__001__4(),
    function ActionValue#(Struct46) rdResp_infoRam__001__3(),
    function ActionValue#(Struct46) rdResp_infoRam__001__2(),
    function ActionValue#(Struct46) rdResp_infoRam__001__1(),
    function ActionValue#(Struct46) rdResp_infoRam__001__0(),
    function Action enq_cp_2__001(Struct45 _),
    function ActionValue#(Struct44) deq_cp_1__001(),
    function Action repGetRq__001(Bit#(9) _),
    function Action rdReq_edirRam__001__3(Bit#(9) _),
    function Action rdReq_edirRam__001__2(Bit#(9) _),
    function Action rdReq_edirRam__001__1(Bit#(9) _),
    function Action rdReq_edirRam__001__0(Bit#(9) _),
    function Action rdReq_infoRam__001__7(Bit#(9) _),
    function Action rdReq_infoRam__001__6(Bit#(9) _),
    function Action rdReq_infoRam__001__5(Bit#(9) _),
    function Action rdReq_infoRam__001__4(Bit#(9) _),
    function Action rdReq_infoRam__001__3(Bit#(9) _),
    function Action rdReq_infoRam__001__2(Bit#(9) _),
    function Action rdReq_infoRam__001__1(Bit#(9) _),
    function Action rdReq_infoRam__001__0(Bit#(9) _),
    function Action enq_cp_1__001(Struct44 _))
    (Module184);
    Reg#(Vector#(4, Struct23)) victims__001 <- mkReg(unpack(0));

    // No rules in this module

    method Action cache__001__infoRq (Bit#(64) x_0);
        let x_1 = (victims__001);
        Struct23 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            let x_3 <- enq_cp_1__001(Struct44 {tag : (x_0)[63:14], index :
            (x_0)[13:5], victim_found : Struct26 {valid : (Bool)'(True), data
            : (Bit#(1))'(1'h0)}});
        end else begin
            Struct23 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                let x_5 <- enq_cp_1__001(Struct44 {tag : (x_0)[63:14], index
                : (x_0)[13:5], victim_found : Struct26 {valid :
                (Bool)'(True), data : (Bit#(1))'(1'h1)}});
            end else begin
                Struct23 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    let x_7 <- enq_cp_1__001(Struct44 {tag : (x_0)[63:14],
                    index : (x_0)[13:5], victim_found : Struct26 {valid :
                    (Bool)'(True), data : (Bit#(1))'(1'h0)}});
                end else begin
                    Struct23 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        let x_9 <- enq_cp_1__001(Struct44 {tag :
                        (x_0)[63:14], index : (x_0)[13:5], victim_found :
                        Struct26 {valid : (Bool)'(True), data :
                        (Bit#(1))'(1'h1)}});
                    end else begin
                        Bit#(9) x_10 = ((x_0)[13:5]);
                        let x_11 <- rdReq_infoRam__001__0(x_10);
                        let x_12 <- rdReq_infoRam__001__1(x_10);
                        let x_13 <- rdReq_infoRam__001__2(x_10);
                        let x_14 <- rdReq_infoRam__001__3(x_10);
                        let x_15 <- rdReq_infoRam__001__4(x_10);
                        let x_16 <- rdReq_infoRam__001__5(x_10);
                        let x_17 <- rdReq_infoRam__001__6(x_10);
                        let x_18 <- rdReq_infoRam__001__7(x_10);
                        let x_19 <- rdReq_edirRam__001__0(x_10);
                        let x_20 <- rdReq_edirRam__001__1(x_10);
                        let x_21 <- rdReq_edirRam__001__2(x_10);
                        let x_22 <- rdReq_edirRam__001__3(x_10);
                        let x_23 <- repGetRq__001(x_10);
                        let x_24 <- enq_cp_1__001(Struct44 {tag :
                        (x_0)[63:14], index : (x_0)[13:5], victim_found :
                        Struct26 {valid : (Bool)'(False), data :
                        unpack(0)}});
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Struct40) cache__001__infoRsValueRq ();
        let x_1 <- deq_cp_1__001();
        Bit#(50) x_2 = ((x_1).tag);
        Bit#(9) x_3 =
        ((x_1).index);
        let x_64 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_4 = (((x_1).victim_found).data);
            let x_5 = (victims__001);
            Struct23 x_6 = ((x_5)[x_4]);
            Struct40 x_7 = (Struct40 {info_index : x_3, info_hit :
            (Bool)'(True), info_way : unpack(0), edir_hit : (Bool)'(False),
            edir_way : unpack(0), edir_slot : Struct41 {valid :
            (Bool)'(False), data : unpack(0)}, info : (x_6).victim_info});
            let x_8 <- enq_cp_2__001(Struct45 {victim_found :
            (x_1).victim_found, may_victim : unpack(0), reps :
            unpack(0)});
            x_64 = x_7;
        end else begin
            Vector#(8, Struct46) x_9 = (unpack(0));
            let x_10 <- rdResp_infoRam__001__0();
            Vector#(8, Struct46) x_11 = (update (x_9, (Bit#(3))'(3'h0),
            x_10));
            let x_12 <- rdResp_infoRam__001__1();
            Vector#(8, Struct46) x_13 = (update (x_11, (Bit#(3))'(3'h1),
            x_12));
            let x_14 <- rdResp_infoRam__001__2();
            Vector#(8, Struct46) x_15 = (update (x_13, (Bit#(3))'(3'h2),
            x_14));
            let x_16 <- rdResp_infoRam__001__3();
            Vector#(8, Struct46) x_17 = (update (x_15, (Bit#(3))'(3'h3),
            x_16));
            let x_18 <- rdResp_infoRam__001__4();
            Vector#(8, Struct46) x_19 = (update (x_17, (Bit#(3))'(3'h4),
            x_18));
            let x_20 <- rdResp_infoRam__001__5();
            Vector#(8, Struct46) x_21 = (update (x_19, (Bit#(3))'(3'h5),
            x_20));
            let x_22 <- rdResp_infoRam__001__6();
            Vector#(8, Struct46) x_23 = (update (x_21, (Bit#(3))'(3'h6),
            x_22));
            let x_24 <- rdResp_infoRam__001__7();
            Vector#(8, Struct46) x_25 = (update (x_23, (Bit#(3))'(3'h7),
            x_24));
            Struct47 x_26 = (((((x_25)[(Bit#(3))'(3'h0)]).tag) == (x_2) ?
            (Struct47 {tm_hit : (Bool)'(True), tm_way : (Bit#(3))'(3'h0),
            tm_value : ((x_25)[(Bit#(3))'(3'h0)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h1)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h1), tm_value :
            ((x_25)[(Bit#(3))'(3'h1)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h2)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h2), tm_value :
            ((x_25)[(Bit#(3))'(3'h2)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h3)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h3), tm_value :
            ((x_25)[(Bit#(3))'(3'h3)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h4)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h4), tm_value :
            ((x_25)[(Bit#(3))'(3'h4)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h5)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h5), tm_value :
            ((x_25)[(Bit#(3))'(3'h5)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h6)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h6), tm_value :
            ((x_25)[(Bit#(3))'(3'h6)]).value}) :
            (((((x_25)[(Bit#(3))'(3'h7)]).tag) == (x_2) ? (Struct47 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(3))'(3'h7), tm_value :
            ((x_25)[(Bit#(3))'(3'h7)]).value}) :
            (unpack(0))))))))))))))))));
            Vector#(4, Struct48) x_27 = (unpack(0));
            let x_28 <- rdResp_edirRam__001__0();
            Vector#(4, Struct48) x_29 = (update (x_27, (Bit#(2))'(2'h0),
            x_28));
            let x_30 <- rdResp_edirRam__001__1();
            Vector#(4, Struct48) x_31 = (update (x_29, (Bit#(2))'(2'h1),
            x_30));
            let x_32 <- rdResp_edirRam__001__2();
            Vector#(4, Struct48) x_33 = (update (x_31, (Bit#(2))'(2'h2),
            x_32));
            let x_34 <- rdResp_edirRam__001__3();
            Vector#(4, Struct48) x_35 = (update (x_33, (Bit#(2))'(2'h3),
            x_34));
            Struct49 x_36 = (((((x_35)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
            (Struct49 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
            tm_value : ((x_35)[(Bit#(2))'(2'h0)]).value}) :
            (((((x_35)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct49 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
            ((x_35)[(Bit#(2))'(2'h1)]).value}) :
            (((((x_35)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct49 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
            ((x_35)[(Bit#(2))'(2'h2)]).value}) :
            (((((x_35)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct49 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
            ((x_35)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
            Struct32 x_37 = ((x_36).tm_value);
            Struct41 x_38 =
            (((((((x_35)[(Bit#(2))'(2'h0)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h0)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h0)}) :
            (((((((x_35)[(Bit#(2))'(2'h1)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h1)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h1)}) :
            (((((((x_35)[(Bit#(2))'(2'h2)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h2)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h2)}) :
            (((((((x_35)[(Bit#(2))'(2'h3)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h0))) ||
            (((((x_35)[(Bit#(2))'(2'h3)]).value).mesi_edir_st) ==
            ((Bit#(3))'(3'h1))) ? (Struct41 {valid : (Bool)'(True), data :
            (Bit#(2))'(2'h3)}) : (Struct41 {valid : (Bool)'(False), data :
            unpack(0)})))))))));
            let x_39 <- repGetRs__001();
            Bit#(3) x_40 = (unpack(0));
            Bit#(8) x_41 = (unpack(0));
            Bit#(3) x_42 = ((! (((x_39)[(Bit#(3))'(3'h7)]) < (x_41)) ?
            ((Bit#(3))'(3'h7)) : (x_40)));
            Bit#(8) x_43 = ((! (((x_39)[(Bit#(3))'(3'h7)]) < (x_41)) ?
            ((x_39)[(Bit#(3))'(3'h7)]) : (x_41)));
            Bit#(3) x_44 = ((! (((x_39)[(Bit#(3))'(3'h6)]) < (x_43)) ?
            ((Bit#(3))'(3'h6)) : (x_42)));
            Bit#(8) x_45 = ((! (((x_39)[(Bit#(3))'(3'h6)]) < (x_43)) ?
            ((x_39)[(Bit#(3))'(3'h6)]) : (x_43)));
            Bit#(3) x_46 = ((! (((x_39)[(Bit#(3))'(3'h5)]) < (x_45)) ?
            ((Bit#(3))'(3'h5)) : (x_44)));
            Bit#(8) x_47 = ((! (((x_39)[(Bit#(3))'(3'h5)]) < (x_45)) ?
            ((x_39)[(Bit#(3))'(3'h5)]) : (x_45)));
            Bit#(3) x_48 = ((! (((x_39)[(Bit#(3))'(3'h4)]) < (x_47)) ?
            ((Bit#(3))'(3'h4)) : (x_46)));
            Bit#(8) x_49 = ((! (((x_39)[(Bit#(3))'(3'h4)]) < (x_47)) ?
            ((x_39)[(Bit#(3))'(3'h4)]) : (x_47)));
            Bit#(3) x_50 = ((! (((x_39)[(Bit#(3))'(3'h3)]) < (x_49)) ?
            ((Bit#(3))'(3'h3)) : (x_48)));
            Bit#(8) x_51 = ((! (((x_39)[(Bit#(3))'(3'h3)]) < (x_49)) ?
            ((x_39)[(Bit#(3))'(3'h3)]) : (x_49)));
            Bit#(3) x_52 = ((! (((x_39)[(Bit#(3))'(3'h2)]) < (x_51)) ?
            ((Bit#(3))'(3'h2)) : (x_50)));
            Bit#(8) x_53 = ((! (((x_39)[(Bit#(3))'(3'h2)]) < (x_51)) ?
            ((x_39)[(Bit#(3))'(3'h2)]) : (x_51)));
            Bit#(3) x_54 = ((! (((x_39)[(Bit#(3))'(3'h1)]) < (x_53)) ?
            ((Bit#(3))'(3'h1)) : (x_52)));
            Bit#(8) x_55 = ((! (((x_39)[(Bit#(3))'(3'h1)]) < (x_53)) ?
            ((x_39)[(Bit#(3))'(3'h1)]) : (x_53)));
            Bit#(3) x_56 = ((! (((x_39)[(Bit#(3))'(3'h0)]) < (x_55)) ?
            ((Bit#(3))'(3'h0)) : (x_54)));
            Bit#(8) x_57 = ((! (((x_39)[(Bit#(3))'(3'h0)]) < (x_55)) ?
            ((x_39)[(Bit#(3))'(3'h0)]) : (x_55)));
            Struct40 x_58 = (Struct40 {info_index : x_3, info_hit :
            (x_26).tm_hit, info_way : (x_26).tm_way, edir_hit :
            (x_36).tm_hit, edir_way : (x_36).tm_way, edir_slot : x_38, info :
            ((x_26).tm_hit ? ((x_26).tm_value) : (Struct11 {mesi_owned :
            (Bool)'(False), mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
            (x_37).mesi_edir_st, mesi_dir_sharers :
            (x_37).mesi_edir_sharers}))});
            Struct46 x_59 = ((x_25)[x_56]);
            Bit#(50) x_60 = ((x_59).tag);
            Struct11 x_61 = ((x_59).value);
            let x_62 <- enq_cp_2__001(Struct45 {victim_found : Struct26
            {valid : (Bool)'(False), data : unpack(0)}, may_victim : Struct28
            {mv_addr : {(x_60),({(x_3),((Bit#(5))'(5'h0))})}, mv_info :
            x_61}, reps : x_39});
            let x_63 <- rdReq_dataRam__001({(((x_26).tm_hit ? ((x_26).tm_way)
            : (x_56))),(x_3)});
            x_64 = x_58;
        end
        return x_64;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__001__valueRsLineRq
    (Struct43 x_0);
        let x_1 <- deq_cp_2__001();
        let x_2 =
        (victims__001);
        let x_61 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_3 = (((x_1).victim_found).data);
            Struct23 x_4 = ((x_2)[x_3]);
            Struct23 x_5 = (Struct23 {victim_valid : (Bool)'(True),
            victim_addr : (x_4).victim_addr, victim_info : ((x_0).info_write
            ? ((x_0).info) : ((x_4).victim_info)), victim_value :
            ((x_0).value_write ? ((x_0).value) : ((x_4).victim_value)),
            victim_req : (x_4).victim_req});
            victims__001 <= update (x_2, x_3, x_5);
            x_61 = (x_4).victim_value;
        end else begin
            let x_6 <- rdResp_dataRam__001();
            Bit#(64) x_7 = ((x_0).addr);
            Bit#(9) x_8 = ((x_7)[13:5]);
            Bit#(3) x_9 = ((x_0).info_way);
            Struct11 x_10 = ((x_0).info);
            Bool x_11 = ((! ((x_10).mesi_owned)) && (((x_10).mesi_status) ==
            ((Bit#(3))'(3'h1))));
            if ((((x_0).info_hit) || (! (x_11))) || ((! ((x_0).edir_hit)) &&
                (x_11)))
                begin
                if ((x_0).info_write) begin
                    Struct50 x_12 = (Struct50 {addr : x_8, datain : Struct46
                    {tag : (x_7)[63:14], value :
                    x_10}});
                    if ((x_9) == ((Bit#(3))'(3'h0))) begin
                        let x_13 <- wrReq_infoRam__001__0(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h1))) begin
                        let x_15 <- wrReq_infoRam__001__1(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h2))) begin
                        let x_17 <- wrReq_infoRam__001__2(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h3))) begin
                        let x_19 <- wrReq_infoRam__001__3(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h4))) begin
                        let x_21 <- wrReq_infoRam__001__4(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h5))) begin
                        let x_23 <- wrReq_infoRam__001__5(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h6))) begin
                        let x_25 <- wrReq_infoRam__001__6(x_12);
                    end else begin

                    end
                    if ((x_9) == ((Bit#(3))'(3'h7))) begin
                        let x_27 <- wrReq_infoRam__001__7(x_12);
                    end else begin

                    end
                    Struct28 x_29 = ((x_1).may_victim);
                    Struct26 x_30 = ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid
                    ? ((((x_2)[(Bit#(1))'(1'h0)]).victim_valid ?
                    ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid ? (Struct26
                    {valid : (Bool)'(False), data : unpack(0)}) : (Struct26
                    {valid : (Bool)'(True), data : (Bit#(1))'(1'h1)}))) :
                    (Struct26 {valid : (Bool)'(True), data :
                    (Bit#(1))'(1'h0)}))) : (Struct26 {valid : (Bool)'(True),
                    data : (Bit#(1))'(1'h1)})));
                    Bit#(1) x_31 = ((x_30).data);
                    victims__001 <= update (x_2, x_31, Struct23 {victim_valid
                    : (Bool)'(True), victim_addr : (x_29).mv_addr,
                    victim_info : (x_29).mv_info, victim_value : x_6,
                    victim_req : Struct14 {valid : (Bool)'(False), data :
                    unpack(0)}});
                    let x_32 <- repAccess__001(Struct51 {acc_type :
                    ((((x_10).mesi_dir_st) == ((Bit#(3))'(3'h0))) ||
                    (((x_10).mesi_dir_st) == ((Bit#(3))'(3'h1))) ?
                    ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))), acc_reps :
                    (x_1).reps, acc_index : x_8, acc_way : x_9});
                end else begin

                end
                if ((x_0).value_write) begin
                    Struct52 x_34 = (Struct52 {addr : {(x_9),((x_7)[13:5])},
                    datain : (x_0).value});
                    let x_35 <- wrReq_dataRam__001(x_34);
                end else begin

                end
            end else begin

            end
            if (((x_0).info_write) && ((x_0).edir_hit)) begin
                Bit#(2) x_38 = ((x_0).edir_way);
                Struct53 x_39 = (Struct53 {addr : (x_7)[13:5], datain :
                Struct48 {tag : (x_7)[63:14], value : (x_11 ? (Struct32
                {mesi_edir_st : (x_10).mesi_dir_st, mesi_edir_sharers :
                (x_10).mesi_dir_sharers}) :
                (unpack(0)))}});
                if ((x_38) == ((Bit#(2))'(2'h0))) begin
                    let x_40 <- wrReq_edirRam__001__0(x_39);
                end else begin

                end
                if ((x_38) == ((Bit#(2))'(2'h1))) begin
                    let x_42 <- wrReq_edirRam__001__1(x_39);
                end else begin

                end
                if ((x_38) == ((Bit#(2))'(2'h2))) begin
                    let x_44 <- wrReq_edirRam__001__2(x_39);
                end else begin

                end
                if ((x_38) == ((Bit#(2))'(2'h3))) begin
                    let x_46 <- wrReq_edirRam__001__3(x_39);
                end else begin

                end
            end else begin
                Struct41 x_48 =
                ((x_0).edir_slot);
                if (((! ((x_0).edir_hit)) && ((x_48).valid)) && (x_11))
                    begin
                    Bit#(2) x_49 = ((x_48).data);
                    Struct53 x_50 = (Struct53 {addr : (x_7)[13:5], datain :
                    Struct48 {tag : (x_7)[63:14], value : Struct32
                    {mesi_edir_st : (x_10).mesi_dir_st, mesi_edir_sharers :
                    (x_10).mesi_dir_sharers}}});
                    if ((x_49) == ((Bit#(2))'(2'h0))) begin
                        let x_51 <- wrReq_edirRam__001__0(x_50);
                    end else begin

                    end
                    if ((x_49) == ((Bit#(2))'(2'h1))) begin
                        let x_53 <- wrReq_edirRam__001__1(x_50);
                    end else begin

                    end
                    if ((x_49) == ((Bit#(2))'(2'h2))) begin
                        let x_55 <- wrReq_edirRam__001__2(x_50);
                    end else begin

                    end
                    if ((x_49) == ((Bit#(2))'(2'h3))) begin
                        let x_57 <- wrReq_edirRam__001__3(x_50);
                    end else begin

                    end
                end else begin

                end
            end
            x_61 = x_6;
        end
        return x_61;
    endmethod

    method ActionValue#(Struct23) cache__001__getVictim ();
        let x_1 = (victims__001);
        Struct38 x_2 = (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        (((((x_1)[(Bit#(1))'(1'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct38 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) : (Struct38 {valid :
        (Bool)'(False), data : unpack(0)})))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method Action cache__001__setVictimRq (Struct24 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(4) x_2 = ((x_0).victim_req);
        let x_3 = (victims__001);
        Struct23 x_4 =
        ((x_3)[(Bit#(1))'(1'h1)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct23 x_5 = (Struct23 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct14 {valid :
            (Bool)'(True), data : x_2}});
            victims__001 <= update (x_3, (Bit#(1))'(1'h1), x_5);
        end else begin
            Struct23 x_6 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct23 x_7 = (Struct23 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct14 {valid : (Bool)'(True), data :
                x_2}});
                victims__001 <= update (x_3, (Bit#(1))'(1'h0), x_7);
            end else begin
                Struct23 x_8 =
                ((x_3)[(Bit#(1))'(1'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct23 x_9 = (Struct23 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct14 {valid :
                    (Bool)'(True), data : x_2}});
                    victims__001 <= update (x_3, (Bit#(1))'(1'h1), x_9);
                end else begin

                end
            end
        end
    endmethod

    method ActionValue#(Bit#(4)) cache__001__releaseVictim (Bit#(64) x_0);
        let x_1 = (victims__001);
        Struct23 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victims__001 <= update (x_1, (Bit#(1))'(1'h0), unpack(0));
            Bit#(4) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct23 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victims__001 <= update (x_1, (Bit#(1))'(1'h1),
                unpack(0));
                Bit#(4) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct23 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victims__001 <= update (x_1, (Bit#(1))'(1'h0),
                    unpack(0));
                    Bit#(4) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct23 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victims__001 <= update (x_1, (Bit#(1))'(1'h1),
                        unpack(0));
                        Bit#(4) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod

    method ActionValue#(Bit#(1)) cache__001__getVictimCount ();
        let x_1 = (victims__001);
        Bit#(1) x_2 = ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((((((x_1)[(Bit#(1))'(1'h0)]).victim_valid)
        && (! ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0)))) +
        ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((Bit#(1))'(1'h0)))));
        return x_2;
    endmethod
endmodule

interface Module185;
    method Action cache__0010__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct60) cache__0010__infoRsValueRq ();
    method ActionValue#(Vector#(4, Bit#(64))) cache__0010__valueRsLineRq
    (Struct64 x_0);
    method ActionValue#(Struct66) cache__0010__getVictim ();
    method Action cache__0010__setVictimRq (Struct67 x_0);
    method ActionValue#(Bit#(3)) cache__0010__releaseVictim (Bit#(64) x_0);
    method ActionValue#(Bit#(1)) cache__0010__getVictimCount ();
endinterface

module mkModule185#(function Action repAccess__0010(Struct74 _),
    function Action wrReq_dataRam__0010(Struct73 _),
    function Action wrReq_infoRam__0010__3(Struct72 _),
    function Action wrReq_infoRam__0010__2(Struct72 _),
    function Action wrReq_infoRam__0010__1(Struct72 _),
    function Action wrReq_infoRam__0010__0(Struct72 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0010(),
    function ActionValue#(Struct69) deq_cp_2__0010(),
    function Action rdReq_dataRam__0010(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__0010(),
    function ActionValue#(Struct70) rdResp_infoRam__0010__3(),
    function ActionValue#(Struct70) rdResp_infoRam__0010__2(),
    function ActionValue#(Struct70) rdResp_infoRam__0010__1(),
    function ActionValue#(Struct70) rdResp_infoRam__0010__0(),
    function Action enq_cp_2__0010(Struct69 _),
    function ActionValue#(Struct68) deq_cp_1__0010(),
    function Action repGetRq__0010(Bit#(8) _),
    function Action rdReq_infoRam__0010__3(Bit#(8) _),
    function Action rdReq_infoRam__0010__2(Bit#(8) _),
    function Action rdReq_infoRam__0010__1(Bit#(8) _),
    function Action rdReq_infoRam__0010__0(Bit#(8) _),
    function Action enq_cp_1__0010(Struct68 _))
    (Module185);
    Reg#(Vector#(4, Struct66)) victims__0010 <- mkReg(unpack(0));

    // No rules in this module

    method Action cache__0010__infoRq (Bit#(64) x_0);
        let x_1 = (victims__0010);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            let x_3 <- enq_cp_1__0010(Struct68 {tag : (x_0)[63:13], index :
            (x_0)[12:5], victim_found : Struct26 {valid : (Bool)'(True), data
            : (Bit#(1))'(1'h0)}});
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                let x_5 <- enq_cp_1__0010(Struct68 {tag : (x_0)[63:13], index
                : (x_0)[12:5], victim_found : Struct26 {valid :
                (Bool)'(True), data : (Bit#(1))'(1'h1)}});
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    let x_7 <- enq_cp_1__0010(Struct68 {tag : (x_0)[63:13],
                    index : (x_0)[12:5], victim_found : Struct26 {valid :
                    (Bool)'(True), data : (Bit#(1))'(1'h0)}});
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        let x_9 <- enq_cp_1__0010(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(True), data :
                        (Bit#(1))'(1'h1)}});
                    end else begin
                        Bit#(8) x_10 = ((x_0)[12:5]);
                        let x_11 <- rdReq_infoRam__0010__0(x_10);
                        let x_12 <- rdReq_infoRam__0010__1(x_10);
                        let x_13 <- rdReq_infoRam__0010__2(x_10);
                        let x_14 <- rdReq_infoRam__0010__3(x_10);
                        let x_15 <- repGetRq__0010(x_10);
                        let x_16 <- enq_cp_1__0010(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(False), data :
                        unpack(0)}});
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Struct60) cache__0010__infoRsValueRq ();
        let x_1 <- deq_cp_1__0010();
        Bit#(51) x_2 = ((x_1).tag);
        Bit#(8) x_3 =
        ((x_1).index);
        let x_36 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_4 = (((x_1).victim_found).data);
            let x_5 = (victims__0010);
            Struct66 x_6 = ((x_5)[x_4]);
            Struct60 x_7 = (Struct60 {info_index : x_3, info_hit :
            (Bool)'(True), info_way : unpack(0), edir_hit : (Bool)'(False),
            edir_way : unpack(0), edir_slot : Struct61 {valid :
            (Bool)'(False), data : unpack(0)}, info : (x_6).victim_info});
            let x_8 <- enq_cp_2__0010(Struct69 {victim_found :
            (x_1).victim_found, may_victim : unpack(0), reps :
            unpack(0)});
            x_36 = x_7;
        end else begin
            Vector#(4, Struct70) x_9 = (unpack(0));
            let x_10 <- rdResp_infoRam__0010__0();
            Vector#(4, Struct70) x_11 = (update (x_9, (Bit#(2))'(2'h0),
            x_10));
            let x_12 <- rdResp_infoRam__0010__1();
            Vector#(4, Struct70) x_13 = (update (x_11, (Bit#(2))'(2'h1),
            x_12));
            let x_14 <- rdResp_infoRam__0010__2();
            Vector#(4, Struct70) x_15 = (update (x_13, (Bit#(2))'(2'h2),
            x_14));
            let x_16 <- rdResp_infoRam__0010__3();
            Vector#(4, Struct70) x_17 = (update (x_15, (Bit#(2))'(2'h3),
            x_16));
            Struct71 x_18 = (((((x_17)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
            (Struct71 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
            tm_value : ((x_17)[(Bit#(2))'(2'h0)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
            ((x_17)[(Bit#(2))'(2'h1)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
            ((x_17)[(Bit#(2))'(2'h2)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
            ((x_17)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
            let x_19 <- repGetRs__0010();
            Bit#(2) x_20 = (unpack(0));
            Bit#(8) x_21 = (unpack(0));
            Bit#(2) x_22 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((Bit#(2))'(2'h3)) : (x_20)));
            Bit#(8) x_23 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((x_19)[(Bit#(2))'(2'h3)]) : (x_21)));
            Bit#(2) x_24 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((Bit#(2))'(2'h2)) : (x_22)));
            Bit#(8) x_25 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((x_19)[(Bit#(2))'(2'h2)]) : (x_23)));
            Bit#(2) x_26 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((Bit#(2))'(2'h1)) : (x_24)));
            Bit#(8) x_27 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((x_19)[(Bit#(2))'(2'h1)]) : (x_25)));
            Bit#(2) x_28 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((Bit#(2))'(2'h0)) : (x_26)));
            Bit#(8) x_29 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((x_19)[(Bit#(2))'(2'h0)]) : (x_27)));
            Struct60 x_30 = (Struct60 {info_index : x_3, info_hit :
            (x_18).tm_hit, info_way : (x_18).tm_way, edir_hit : unpack(0),
            edir_way : unpack(0), edir_slot : unpack(0), info :
            (x_18).tm_value});
            Struct70 x_31 = ((x_17)[x_28]);
            Bit#(51) x_32 = ((x_31).tag);
            Struct11 x_33 = ((x_31).value);
            let x_34 <- enq_cp_2__0010(Struct69 {victim_found : Struct26
            {valid : (Bool)'(False), data : unpack(0)}, may_victim : Struct28
            {mv_addr : {(x_32),({(x_3),((Bit#(5))'(5'h0))})}, mv_info :
            x_33}, reps : x_19});
            let x_35 <- rdReq_dataRam__0010({(((x_18).tm_hit ?
            ((x_18).tm_way) : (x_28))),(x_3)});
            x_36 = x_30;
        end
        return x_36;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__0010__valueRsLineRq
    (Struct64 x_0);
        let x_1 <- deq_cp_2__0010();
        let x_2 =
        (victims__0010);
        let x_29 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_3 = (((x_1).victim_found).data);
            Struct66 x_4 = ((x_2)[x_3]);
            Struct66 x_5 = (Struct66 {victim_valid : (Bool)'(True),
            victim_addr : (x_4).victim_addr, victim_info : ((x_0).info_write
            ? ((x_0).info) : ((x_4).victim_info)), victim_value :
            ((x_0).value_write ? ((x_0).value) : ((x_4).victim_value)),
            victim_req : (x_4).victim_req});
            victims__0010 <= update (x_2, x_3, x_5);
            x_29 = (x_4).victim_value;
        end else begin
            let x_6 <- rdResp_dataRam__0010();
            Bit#(64) x_7 = ((x_0).addr);
            Bit#(8) x_8 = ((x_7)[12:5]);
            Bit#(2) x_9 = ((x_0).info_way);
            Struct11 x_10 =
            ((x_0).info);
            if ((x_0).info_write) begin
                Struct72 x_11 = (Struct72 {addr : x_8, datain : Struct70 {tag
                : (x_7)[63:13], value :
                x_10}});
                if ((x_9) == ((Bit#(2))'(2'h0))) begin
                    let x_12 <- wrReq_infoRam__0010__0(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h1))) begin
                    let x_14 <- wrReq_infoRam__0010__1(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h2))) begin
                    let x_16 <- wrReq_infoRam__0010__2(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h3))) begin
                    let x_18 <- wrReq_infoRam__0010__3(x_11);
                end else begin

                end
                if ((x_0).value_write) begin
                    Struct73 x_20 = (Struct73 {addr : {(x_9),((x_7)[12:5])},
                    datain : (x_0).value});
                    let x_21 <- wrReq_dataRam__0010(x_20);
                end else begin

                end
                if (! ((x_0).info_hit)) begin
                    Struct28 x_23 = ((x_1).may_victim);
                    Struct26 x_24 = ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid
                    ? ((((x_2)[(Bit#(1))'(1'h0)]).victim_valid ?
                    ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid ? (Struct26
                    {valid : (Bool)'(False), data : unpack(0)}) : (Struct26
                    {valid : (Bool)'(True), data : (Bit#(1))'(1'h1)}))) :
                    (Struct26 {valid : (Bool)'(True), data :
                    (Bit#(1))'(1'h0)}))) : (Struct26 {valid : (Bool)'(True),
                    data : (Bit#(1))'(1'h1)})));
                    Bit#(1) x_25 = ((x_24).data);
                    victims__0010 <= update (x_2, x_25, Struct66
                    {victim_valid : (Bool)'(True), victim_addr :
                    (x_23).mv_addr, victim_info : (x_23).mv_info,
                    victim_value : x_6, victim_req : Struct10 {valid :
                    (Bool)'(False), data : unpack(0)}});
                end else begin

                end
                let x_27 <- repAccess__0010(Struct74 {acc_type :
                ((((x_10).mesi_dir_st) == ((Bit#(3))'(3'h0))) ||
                (((x_10).mesi_dir_st) == ((Bit#(3))'(3'h1))) ?
                ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))), acc_reps :
                (x_1).reps, acc_index : x_8, acc_way : x_9});
            end else begin

            end
            x_29 = x_6;
        end
        return x_29;
    endmethod

    method ActionValue#(Struct66) cache__0010__getVictim ();
        let x_1 = (victims__0010);
        Struct75 x_2 = (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        (((((x_1)[(Bit#(1))'(1'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) : (Struct75 {valid :
        (Bool)'(False), data : unpack(0)})))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method Action cache__0010__setVictimRq (Struct67 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victims__0010);
        Struct66 x_4 =
        ((x_3)[(Bit#(1))'(1'h1)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct66 x_5 = (Struct66 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct10 {valid :
            (Bool)'(True), data : x_2}});
            victims__0010 <= update (x_3, (Bit#(1))'(1'h1), x_5);
        end else begin
            Struct66 x_6 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct66 x_7 = (Struct66 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct10 {valid : (Bool)'(True), data :
                x_2}});
                victims__0010 <= update (x_3, (Bit#(1))'(1'h0), x_7);
            end else begin
                Struct66 x_8 =
                ((x_3)[(Bit#(1))'(1'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct66 x_9 = (Struct66 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct10 {valid :
                    (Bool)'(True), data : x_2}});
                    victims__0010 <= update (x_3, (Bit#(1))'(1'h1), x_9);
                end else begin

                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) cache__0010__releaseVictim (Bit#(64) x_0);
        let x_1 = (victims__0010);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victims__0010 <= update (x_1, (Bit#(1))'(1'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victims__0010 <= update (x_1, (Bit#(1))'(1'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victims__0010 <= update (x_1, (Bit#(1))'(1'h0),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victims__0010 <= update (x_1, (Bit#(1))'(1'h1),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod

    method ActionValue#(Bit#(1)) cache__0010__getVictimCount ();
        let x_1 = (victims__0010);
        Bit#(1) x_2 = ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((((((x_1)[(Bit#(1))'(1'h0)]).victim_valid)
        && (! ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0)))) +
        ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((Bit#(1))'(1'h0)))));
        return x_2;
    endmethod
endmodule

interface Module186;
    method Action cache__0011__infoRq (Bit#(64) x_0);
    method ActionValue#(Struct60) cache__0011__infoRsValueRq ();
    method ActionValue#(Vector#(4, Bit#(64))) cache__0011__valueRsLineRq
    (Struct64 x_0);
    method ActionValue#(Struct66) cache__0011__getVictim ();
    method Action cache__0011__setVictimRq (Struct67 x_0);
    method ActionValue#(Bit#(3)) cache__0011__releaseVictim (Bit#(64) x_0);
    method ActionValue#(Bit#(1)) cache__0011__getVictimCount ();
endinterface

module mkModule186#(function Action repAccess__0011(Struct74 _),
    function Action wrReq_dataRam__0011(Struct73 _),
    function Action wrReq_infoRam__0011__3(Struct72 _),
    function Action wrReq_infoRam__0011__2(Struct72 _),
    function Action wrReq_infoRam__0011__1(Struct72 _),
    function Action wrReq_infoRam__0011__0(Struct72 _),
    function ActionValue#(Vector#(4, Bit#(64))) rdResp_dataRam__0011(),
    function ActionValue#(Struct69) deq_cp_2__0011(),
    function Action rdReq_dataRam__0011(Bit#(10) _),
    function ActionValue#(Vector#(4, Bit#(8))) repGetRs__0011(),
    function ActionValue#(Struct70) rdResp_infoRam__0011__3(),
    function ActionValue#(Struct70) rdResp_infoRam__0011__2(),
    function ActionValue#(Struct70) rdResp_infoRam__0011__1(),
    function ActionValue#(Struct70) rdResp_infoRam__0011__0(),
    function Action enq_cp_2__0011(Struct69 _),
    function ActionValue#(Struct68) deq_cp_1__0011(),
    function Action repGetRq__0011(Bit#(8) _),
    function Action rdReq_infoRam__0011__3(Bit#(8) _),
    function Action rdReq_infoRam__0011__2(Bit#(8) _),
    function Action rdReq_infoRam__0011__1(Bit#(8) _),
    function Action rdReq_infoRam__0011__0(Bit#(8) _),
    function Action enq_cp_1__0011(Struct68 _))
    (Module186);
    Reg#(Vector#(4, Struct66)) victims__0011 <- mkReg(unpack(0));

    // No rules in this module

    method Action cache__0011__infoRq (Bit#(64) x_0);
        let x_1 = (victims__0011);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0))) begin
            let x_3 <- enq_cp_1__0011(Struct68 {tag : (x_0)[63:13], index :
            (x_0)[12:5], victim_found : Struct26 {valid : (Bool)'(True), data
            : (Bit#(1))'(1'h0)}});
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                let x_5 <- enq_cp_1__0011(Struct68 {tag : (x_0)[63:13], index
                : (x_0)[12:5], victim_found : Struct26 {valid :
                (Bool)'(True), data : (Bit#(1))'(1'h1)}});
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    let x_7 <- enq_cp_1__0011(Struct68 {tag : (x_0)[63:13],
                    index : (x_0)[12:5], victim_found : Struct26 {valid :
                    (Bool)'(True), data : (Bit#(1))'(1'h0)}});
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        let x_9 <- enq_cp_1__0011(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(True), data :
                        (Bit#(1))'(1'h1)}});
                    end else begin
                        Bit#(8) x_10 = ((x_0)[12:5]);
                        let x_11 <- rdReq_infoRam__0011__0(x_10);
                        let x_12 <- rdReq_infoRam__0011__1(x_10);
                        let x_13 <- rdReq_infoRam__0011__2(x_10);
                        let x_14 <- rdReq_infoRam__0011__3(x_10);
                        let x_15 <- repGetRq__0011(x_10);
                        let x_16 <- enq_cp_1__0011(Struct68 {tag :
                        (x_0)[63:13], index : (x_0)[12:5], victim_found :
                        Struct26 {valid : (Bool)'(False), data :
                        unpack(0)}});
                    end
                end
            end
        end
    endmethod

    method ActionValue#(Struct60) cache__0011__infoRsValueRq ();
        let x_1 <- deq_cp_1__0011();
        Bit#(51) x_2 = ((x_1).tag);
        Bit#(8) x_3 =
        ((x_1).index);
        let x_36 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_4 = (((x_1).victim_found).data);
            let x_5 = (victims__0011);
            Struct66 x_6 = ((x_5)[x_4]);
            Struct60 x_7 = (Struct60 {info_index : x_3, info_hit :
            (Bool)'(True), info_way : unpack(0), edir_hit : (Bool)'(False),
            edir_way : unpack(0), edir_slot : Struct61 {valid :
            (Bool)'(False), data : unpack(0)}, info : (x_6).victim_info});
            let x_8 <- enq_cp_2__0011(Struct69 {victim_found :
            (x_1).victim_found, may_victim : unpack(0), reps :
            unpack(0)});
            x_36 = x_7;
        end else begin
            Vector#(4, Struct70) x_9 = (unpack(0));
            let x_10 <- rdResp_infoRam__0011__0();
            Vector#(4, Struct70) x_11 = (update (x_9, (Bit#(2))'(2'h0),
            x_10));
            let x_12 <- rdResp_infoRam__0011__1();
            Vector#(4, Struct70) x_13 = (update (x_11, (Bit#(2))'(2'h1),
            x_12));
            let x_14 <- rdResp_infoRam__0011__2();
            Vector#(4, Struct70) x_15 = (update (x_13, (Bit#(2))'(2'h2),
            x_14));
            let x_16 <- rdResp_infoRam__0011__3();
            Vector#(4, Struct70) x_17 = (update (x_15, (Bit#(2))'(2'h3),
            x_16));
            Struct71 x_18 = (((((x_17)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
            (Struct71 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
            tm_value : ((x_17)[(Bit#(2))'(2'h0)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
            ((x_17)[(Bit#(2))'(2'h1)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
            ((x_17)[(Bit#(2))'(2'h2)]).value}) :
            (((((x_17)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct71 {tm_hit :
            (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
            ((x_17)[(Bit#(2))'(2'h3)]).value}) : (unpack(0))))))))));
            let x_19 <- repGetRs__0011();
            Bit#(2) x_20 = (unpack(0));
            Bit#(8) x_21 = (unpack(0));
            Bit#(2) x_22 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((Bit#(2))'(2'h3)) : (x_20)));
            Bit#(8) x_23 = ((! (((x_19)[(Bit#(2))'(2'h3)]) < (x_21)) ?
            ((x_19)[(Bit#(2))'(2'h3)]) : (x_21)));
            Bit#(2) x_24 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((Bit#(2))'(2'h2)) : (x_22)));
            Bit#(8) x_25 = ((! (((x_19)[(Bit#(2))'(2'h2)]) < (x_23)) ?
            ((x_19)[(Bit#(2))'(2'h2)]) : (x_23)));
            Bit#(2) x_26 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((Bit#(2))'(2'h1)) : (x_24)));
            Bit#(8) x_27 = ((! (((x_19)[(Bit#(2))'(2'h1)]) < (x_25)) ?
            ((x_19)[(Bit#(2))'(2'h1)]) : (x_25)));
            Bit#(2) x_28 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((Bit#(2))'(2'h0)) : (x_26)));
            Bit#(8) x_29 = ((! (((x_19)[(Bit#(2))'(2'h0)]) < (x_27)) ?
            ((x_19)[(Bit#(2))'(2'h0)]) : (x_27)));
            Struct60 x_30 = (Struct60 {info_index : x_3, info_hit :
            (x_18).tm_hit, info_way : (x_18).tm_way, edir_hit : unpack(0),
            edir_way : unpack(0), edir_slot : unpack(0), info :
            (x_18).tm_value});
            Struct70 x_31 = ((x_17)[x_28]);
            Bit#(51) x_32 = ((x_31).tag);
            Struct11 x_33 = ((x_31).value);
            let x_34 <- enq_cp_2__0011(Struct69 {victim_found : Struct26
            {valid : (Bool)'(False), data : unpack(0)}, may_victim : Struct28
            {mv_addr : {(x_32),({(x_3),((Bit#(5))'(5'h0))})}, mv_info :
            x_33}, reps : x_19});
            let x_35 <- rdReq_dataRam__0011({(((x_18).tm_hit ?
            ((x_18).tm_way) : (x_28))),(x_3)});
            x_36 = x_30;
        end
        return x_36;
    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) cache__0011__valueRsLineRq
    (Struct64 x_0);
        let x_1 <- deq_cp_2__0011();
        let x_2 =
        (victims__0011);
        let x_29 = ?;
        if (((x_1).victim_found).valid) begin
            Bit#(1) x_3 = (((x_1).victim_found).data);
            Struct66 x_4 = ((x_2)[x_3]);
            Struct66 x_5 = (Struct66 {victim_valid : (Bool)'(True),
            victim_addr : (x_4).victim_addr, victim_info : ((x_0).info_write
            ? ((x_0).info) : ((x_4).victim_info)), victim_value :
            ((x_0).value_write ? ((x_0).value) : ((x_4).victim_value)),
            victim_req : (x_4).victim_req});
            victims__0011 <= update (x_2, x_3, x_5);
            x_29 = (x_4).victim_value;
        end else begin
            let x_6 <- rdResp_dataRam__0011();
            Bit#(64) x_7 = ((x_0).addr);
            Bit#(8) x_8 = ((x_7)[12:5]);
            Bit#(2) x_9 = ((x_0).info_way);
            Struct11 x_10 =
            ((x_0).info);
            if ((x_0).info_write) begin
                Struct72 x_11 = (Struct72 {addr : x_8, datain : Struct70 {tag
                : (x_7)[63:13], value :
                x_10}});
                if ((x_9) == ((Bit#(2))'(2'h0))) begin
                    let x_12 <- wrReq_infoRam__0011__0(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h1))) begin
                    let x_14 <- wrReq_infoRam__0011__1(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h2))) begin
                    let x_16 <- wrReq_infoRam__0011__2(x_11);
                end else begin

                end
                if ((x_9) == ((Bit#(2))'(2'h3))) begin
                    let x_18 <- wrReq_infoRam__0011__3(x_11);
                end else begin

                end
                if ((x_0).value_write) begin
                    Struct73 x_20 = (Struct73 {addr : {(x_9),((x_7)[12:5])},
                    datain : (x_0).value});
                    let x_21 <- wrReq_dataRam__0011(x_20);
                end else begin

                end
                if (! ((x_0).info_hit)) begin
                    Struct28 x_23 = ((x_1).may_victim);
                    Struct26 x_24 = ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid
                    ? ((((x_2)[(Bit#(1))'(1'h0)]).victim_valid ?
                    ((((x_2)[(Bit#(1))'(1'h1)]).victim_valid ? (Struct26
                    {valid : (Bool)'(False), data : unpack(0)}) : (Struct26
                    {valid : (Bool)'(True), data : (Bit#(1))'(1'h1)}))) :
                    (Struct26 {valid : (Bool)'(True), data :
                    (Bit#(1))'(1'h0)}))) : (Struct26 {valid : (Bool)'(True),
                    data : (Bit#(1))'(1'h1)})));
                    Bit#(1) x_25 = ((x_24).data);
                    victims__0011 <= update (x_2, x_25, Struct66
                    {victim_valid : (Bool)'(True), victim_addr :
                    (x_23).mv_addr, victim_info : (x_23).mv_info,
                    victim_value : x_6, victim_req : Struct10 {valid :
                    (Bool)'(False), data : unpack(0)}});
                end else begin

                end
                let x_27 <- repAccess__0011(Struct74 {acc_type :
                ((((x_10).mesi_dir_st) == ((Bit#(3))'(3'h0))) ||
                (((x_10).mesi_dir_st) == ((Bit#(3))'(3'h1))) ?
                ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))), acc_reps :
                (x_1).reps, acc_index : x_8, acc_way : x_9});
            end else begin

            end
            x_29 = x_6;
        end
        return x_29;
    endmethod

    method ActionValue#(Struct66) cache__0011__getVictim ();
        let x_1 = (victims__0011);
        Struct75 x_2 = (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        (((((x_1)[(Bit#(1))'(1'h0)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? (Struct75 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) : (Struct75 {valid :
        (Bool)'(False), data : unpack(0)})))))));
        when ((x_2).valid, noAction);
        return (x_2).data;
    endmethod

    method Action cache__0011__setVictimRq (Struct67 x_0);
        Bit#(64) x_1 = ((x_0).victim_addr);
        Bit#(3) x_2 = ((x_0).victim_req);
        let x_3 = (victims__0011);
        Struct66 x_4 =
        ((x_3)[(Bit#(1))'(1'h1)]);
        if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_1)))
            begin
            Struct66 x_5 = (Struct66 {victim_valid : (x_4).victim_valid,
            victim_addr : (x_4).victim_addr, victim_info : (x_4).victim_info,
            victim_value : (x_4).victim_value, victim_req : Struct10 {valid :
            (Bool)'(True), data : x_2}});
            victims__0011 <= update (x_3, (Bit#(1))'(1'h1), x_5);
        end else begin
            Struct66 x_6 =
            ((x_3)[(Bit#(1))'(1'h0)]);
            if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_1)))
                begin
                Struct66 x_7 = (Struct66 {victim_valid : (x_6).victim_valid,
                victim_addr : (x_6).victim_addr, victim_info :
                (x_6).victim_info, victim_value : (x_6).victim_value,
                victim_req : Struct10 {valid : (Bool)'(True), data :
                x_2}});
                victims__0011 <= update (x_3, (Bit#(1))'(1'h0), x_7);
            end else begin
                Struct66 x_8 =
                ((x_3)[(Bit#(1))'(1'h1)]);
                if (((x_8).victim_valid) && (((x_8).victim_addr) == (x_1)))
                    begin
                    Struct66 x_9 = (Struct66 {victim_valid :
                    (x_8).victim_valid, victim_addr : (x_8).victim_addr,
                    victim_info : (x_8).victim_info, victim_value :
                    (x_8).victim_value, victim_req : Struct10 {valid :
                    (Bool)'(True), data : x_2}});
                    victims__0011 <= update (x_3, (Bit#(1))'(1'h1), x_9);
                end else begin

                end
            end
        end
    endmethod

    method ActionValue#(Bit#(3)) cache__0011__releaseVictim (Bit#(64) x_0);
        let x_1 = (victims__0011);
        Struct66 x_2 =
        ((x_1)[(Bit#(1))'(1'h0)]);
        let x_13 = ?;
        if (((x_2).victim_valid) && (((x_2).victim_addr) == (x_0)))
            begin
            victims__0011 <= update (x_1, (Bit#(1))'(1'h0),
            unpack(0));
            Bit#(3) x_3 = (((x_2).victim_req).data);
            x_13 = x_3;
        end else begin
            Struct66 x_4 =
            ((x_1)[(Bit#(1))'(1'h1)]);
            let x_12 = ?;
            if (((x_4).victim_valid) && (((x_4).victim_addr) == (x_0)))
                begin
                victims__0011 <= update (x_1, (Bit#(1))'(1'h1),
                unpack(0));
                Bit#(3) x_5 = (((x_4).victim_req).data);
                x_12 = x_5;
            end else begin
                Struct66 x_6 =
                ((x_1)[(Bit#(1))'(1'h0)]);
                let x_11 = ?;
                if (((x_6).victim_valid) && (((x_6).victim_addr) == (x_0)))
                    begin
                    victims__0011 <= update (x_1, (Bit#(1))'(1'h0),
                    unpack(0));
                    Bit#(3) x_7 = (((x_6).victim_req).data);
                    x_11 = x_7;
                end else begin
                    Struct66 x_8 =
                    ((x_1)[(Bit#(1))'(1'h1)]);
                    let x_10 = ?;
                    if (((x_8).victim_valid) && (((x_8).victim_addr) ==
                        (x_0))) begin
                        victims__0011 <= update (x_1, (Bit#(1))'(1'h1),
                        unpack(0));
                        Bit#(3) x_9 = (((x_8).victim_req).data);
                        x_10 = x_9;
                    end else begin
                        x_10 = unpack(0);
                    end
                    x_11 = x_10;
                end
                x_12 = x_11;
            end
            x_13 = x_12;
        end
        return x_13;
    endmethod

    method ActionValue#(Bit#(1)) cache__0011__getVictimCount ();
        let x_1 = (victims__0011);
        Bit#(1) x_2 = ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((((((x_1)[(Bit#(1))'(1'h0)]).victim_valid)
        && (! ((((x_1)[(Bit#(1))'(1'h0)]).victim_req).valid)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0)))) +
        ((((((x_1)[(Bit#(1))'(1'h1)]).victim_valid) && (!
        ((((x_1)[(Bit#(1))'(1'h1)]).victim_req).valid)) ? ((Bit#(1))'(1'h1))
        : ((Bit#(1))'(1'h0)))) + ((Bit#(1))'(1'h0)))));
        return x_2;
    endmethod
endmodule

interface Module187;

endinterface

module mkModule187#(function Action cache__00__setVictimRq(Struct24 _),
    function ActionValue#(Bit#(4)) getULImm_00(Struct1 _),
    function ActionValue#(Struct23) cache__00__getVictim(),
    function Action transferUpDown_00(Struct22 _),
    function Action broadcast_parentChildren00(Struct20 _),
    function Action registerDL_00(Struct19 _),
    function Action registerUL_00(Struct18 _),
    function ActionValue#(Bit#(1)) cache__00__getVictimCount(),
    function ActionValue#(Bit#(4)) getULCount_00(),
    function Action makeEnq_parentChildren00(Struct17 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__00__valueRsLineRq(Struct16 _),
    function ActionValue#(Struct13) getMSHR_00(Bit#(4) _),
    function ActionValue#(Struct12) deq_fifoL2E00(),
    function Action enq_fifoL2E00(Struct12 _),
    function ActionValue#(Struct9) cache__00__infoRsValueRq(),
    function ActionValue#(Struct3) deq_fifoI2L00(),
    function ActionValue#(Struct8) getRsReady_00(),
    function Action releaseMSHR_00(Bit#(4) _),
    function ActionValue#(Bit#(4)) cache__00__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct7) getWait_00(),
    function Action addRs_00(Struct6 _),
    function ActionValue#(Struct5) getCRqSlot_00(Struct4 _),
    function ActionValue#(Bit#(4)) findUL_00(Bit#(64) _),
    function Action enq_fifoI2L00(Struct3 _),
    function Action cache__00__infoRq(Bit#(64) _),
    function ActionValue#(Struct5) getPRqSlot_00(Struct4 _),
    function ActionValue#(Struct3) deq_fifoInput00())
    (Module187);

    rule rule_ir_prq_00;
        let x_0 <- deq_fifoInput00();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_00(Struct4 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).ir_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__00__infoRq((x_2).addr);
            Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L00(x_5);
        end else begin

        end
    endrule

    rule rule_ir_prs_00;
        let x_0 <- deq_fifoInput00();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- findUL_00((x_2).addr);
        let x_4 <- cache__00__infoRq((x_2).addr);
        Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : x_3});
        let x_6 <- enq_fifoI2L00(x_5);
    endrule

    rule rule_ir_crq_00;
        let x_0 <- deq_fifoInput00();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getCRqSlot_00(Struct4 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__00__infoRq((x_2).addr);
            Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L00(x_5);
        end else begin

        end
    endrule

    rule rule_ir_crs_00;
        let x_0 <- deq_fifoInput00();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_00(Struct6 {r_dl_midx : (x_1)[0:0], r_dl_msg :
        x_2});
    endrule

    rule rule_ir_retry_00;
        let x_0 <- getWait_00();
        when ((x_0).valid, noAction);
        Struct4 x_1 = ((x_0).data);
        Struct1 x_2 = ((x_1).r_msg);
        let x_3 <- cache__00__infoRq((x_2).addr);
        Struct3 x_4 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg : x_2,
        ir_msg_from : (x_1).r_msg_from, ir_mshr_id : (x_1).r_id});
        let x_5 <- enq_fifoI2L00(x_4);
    endrule

    rule rule_ir_invrs_00;
        let x_0 <- deq_fifoInput00();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- cache__00__releaseVictim((x_2).addr);
        let x_4 <- releaseMSHR_00(x_3);
    endrule

    rule rule_ir_rsrel_00;
        let x_0 <- getRsReady_00();
        Struct1 x_1 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        let x_2 <- cache__00__infoRq((x_0).r_addr);
        Struct3 x_3 = (Struct3 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_1,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id});
        let x_4 <- enq_fifoI2L00(x_3);
    endrule

    rule rule_lr_00;
        let x_0 <- deq_fifoI2L00();
        let x_1 <- cache__00__infoRsValueRq();
        Struct12 x_2 = (Struct12 {lr_ir_pp : x_0, lr_ir : x_1});
        let x_3 <- enq_fifoL2E00(x_2);
    endrule

    rule rule_exec_00_000000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_12).dir_st))) && ((x_11) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) :
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))}).dir_excl)))},
        value_write : (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_16}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_001000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_01000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_00();
        let x_17 <- cache__00__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_00(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
    endrule

    rule rule_exec_00_03000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_10000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) || (((x_11) ==
        ((Bit#(3))'(3'h2))) && (((x_10) == ((Bool)'(True))) &&
        ((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) ==
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        let x_18 <- cache__00__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
    endrule

    rule rule_exec_00_11000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_00();
        let x_17 <- cache__00__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_00(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
    endrule

    rule rule_exec_00_14000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_15000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))) == ((Bit#(2))'(2'h0)))) && (((x_10) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_11))) &&
        (((x_12).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        let x_17 <- broadcast_parentChildren00(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_25000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren00(x_16);
    endrule

    rule rule_exec_00_2600000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_2601000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_261000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_27000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_28000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren00(x_16);
    endrule

    rule rule_exec_00_290000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_291000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_210000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_211000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value});
        let x_19 <- cache__00__valueRsLineRq(x_18);
        Struct17 x_20 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_040000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_070000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_1600000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_1601000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_11000000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_11001000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_11002000;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_000001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_12).dir_st))) && ((x_11) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) :
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))}).dir_excl)))},
        value_write : (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_16}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_001001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_01001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_00();
        let x_17 <- cache__00__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_00(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h5))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
    endrule

    rule rule_exec_00_03001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_10001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) || (((x_11) ==
        ((Bit#(3))'(3'h2))) && (((x_10) == ((Bool)'(True))) &&
        ((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) ==
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        let x_18 <- cache__00__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
    endrule

    rule rule_exec_00_11001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_00();
        let x_17 <- cache__00__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_00(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h5))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
    endrule

    rule rule_exec_00_14001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_15001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))) == ((Bit#(2))'(2'h0)))) && (((x_10) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_11))) &&
        (((x_12).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        let x_17 <- broadcast_parentChildren00(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_25001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren00(x_16);
    endrule

    rule rule_exec_00_2600001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_2601001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_261001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_27001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_28001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren00(x_16);
    endrule

    rule rule_exec_00_290001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_291001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__00__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_210001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_211001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value});
        let x_19 <- cache__00__valueRsLineRq(x_18);
        Struct17 x_20 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
    endrule

    rule rule_exec_00_040001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_070001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_1600001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_1601001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_11000001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_11001001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_11002001;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- addRs_00(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_00_020;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct16 x_16 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_excl)))}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct16 x_19 = (Struct16 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct16 x_20 = (Struct16 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_21 <- cache__00__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_00(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_24 <- makeEnq_parentChildren00(x_23);
    endrule

    rule rule_exec_00_021;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct16 x_16 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct16 x_19 = (Struct16 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct16 x_20 = (Struct16 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_21 <- cache__00__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_00(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_24 <- makeEnq_parentChildren00(x_23);
    endrule

    rule rule_exec_00_041;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct21 x_13 = (Struct21 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_8).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))))}, msg :
        ((x_8).m_dl_rss)[((((x_8).m_dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        (unpack(0)))))))]});
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ((x_8).m_qidx);
        Struct16 x_16 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : ((unpack(0)) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_st, mesi_dir_sharers : (((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        ((unpack(0)) | (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_st) ==
        ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : unpack(0), dir_sharers : ((unpack(0)) | (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0]))) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : ((unpack(0)) | (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_excl)))},
        value_write : (x_16).value_write, value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct16 x_19 = (Struct16 {addr : (x_18).addr, info_write :
        (x_18).info_write, info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : (x_18).info,
        value_write : (Bool)'(True), value : ((x_13).msg).value});
        Struct16 x_20 = (Struct16 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_19).info).mesi_status,
        mesi_dir_st : ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache__00__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_00(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_14).addr, value :
        ((x_13).msg).value}});
        let x_24 <- makeEnq_parentChildren00(x_23);
    endrule

    rule rule_exec_00_05;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_12).dir_st))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_06;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_11))) && ((!
        (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_12).dir_st))))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h2)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_071;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct21 x_13 = (Struct21 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_8).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))))}, msg :
        ((x_8).m_dl_rss)[((((x_8).m_dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        (unpack(0)))))))]});
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ((x_8).m_qidx);
        Struct16 x_16 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : (unpack(0)) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_st,
        mesi_dir_sharers : (((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        unpack(0), dir_sharers : (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct16 x_19 = (Struct16 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct16 x_20 = (Struct16 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : ((x_13).msg).value});
        let x_21 <- cache__00__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_00(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_14).addr, value :
        ((x_13).msg).value}});
        let x_24 <- makeEnq_parentChildren00(x_23);
    endrule

    rule rule_exec_00_12;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((((x_12).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << (({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])})[0:0])))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct16 x_16 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct16 x_19 = (Struct16 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        let x_20 <- cache__00__valueRsLineRq(x_19);
        let x_21 <- releaseMSHR_00(x_4);
        Struct17 x_22 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
    endrule

    rule rule_exec_00_13;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])})[0:0])))) ==
        ((Bit#(2))'(2'h0)))) && (((x_12).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct16 x_15 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_15).info).mesi_status,
        mesi_dir_st : ((x_15).info).mesi_dir_st, mesi_dir_sharers :
        ((x_15).info).mesi_dir_sharers}, value_write : (x_15).value_write,
        value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        let x_18 <- transferUpDown_00(Struct22 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((x_14)[0:0])))});
        let x_19 <- broadcast_parentChildren00(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((x_14)[0:0]))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_161;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct16 x_15 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__00__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_00(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
    endrule

    rule rule_exec_00_170;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_171;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
    endrule

    rule rule_exec_00_190;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (x_12).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(3))'(3'h2)});
        let x_17 <- broadcast_parentChildren00(Struct20 {cs_inds :
        (x_12).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_191;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h2)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
    endrule

    rule rule_exec_00_192;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__00__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_00(Struct19 {r_id : x_4, r_dl_rss_from :
        (x_12).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(3))'(3'h2)});
        let x_17 <- broadcast_parentChildren00(Struct20 {cs_inds :
        (x_12).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_00_11010;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct16 x_15 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__00__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_00(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
    endrule

    rule rule_exec_00_11011;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct16 x_15 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct16 x_17 = (Struct16 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct16 x_18 = (Struct16 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__00__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_00(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
    endrule

    rule rule_exec_00_20;
        let x_0 <- cache__00__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_00(x_4);
        let x_6 <- cache__00__setVictimRq(Struct24 {victim_addr : x_1,
        victim_req : x_5});
        Struct13 x_7 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_9) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_10))
        && ((x_10) < ((Bit#(3))'(3'h4)))) && (((x_11).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        let x_12 <- registerUL_00(Struct18 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_14 <- makeEnq_parentChildren00(x_13);
    endrule

    rule rule_exec_00_21;
        let x_0 <- cache__00__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_00(x_4);
        let x_6 <- cache__00__setVictimRq(Struct24 {victim_addr : x_1,
        victim_req : x_5});
        Struct13 x_7 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when ((((x_11).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_9) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_10))) || (((x_9) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_10)) && ((x_10) <
        ((Bit#(3))'(3'h3)))))), noAction);
        let x_12 <- registerUL_00(Struct18 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_14 <- makeEnq_parentChildren00(x_13);
    endrule

    rule rule_exec_00_22;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h16)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when (! ((x_8).m_rsb), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct16 x_14 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_15 = (Struct16 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct16 x_16 = (Struct16 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__00__valueRsLineRq(x_16);
        let x_18 <- releaseMSHR_00(x_4);
    endrule

    rule rule_exec_00_23;
        let x_0 <- deq_fifoL2E00();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct9 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_00(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((((x_11) == ((Bit#(3))'(3'h1))) && (! (((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_11) == ((Bit#(3))'(3'h2))) && ((x_10)
        == ((Bool)'(False)))), noAction);
        Struct16 x_13 = (Struct16 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct16 x_14 = (Struct16 {addr : (x_13).addr, info_write :
        (Bool)'(True), info_hit : (x_13).info_hit, info_way :
        (x_13).info_way, edir_hit : (x_13).edir_hit, edir_way :
        (x_13).edir_way, edir_slot : (x_13).edir_slot, info : Struct11
        {mesi_owned : ((x_13).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_13).info).mesi_dir_st,
        mesi_dir_sharers : ((x_13).info).mesi_dir_sharers}, value_write :
        (x_13).value_write, value : (x_13).value});
        let x_15 <- cache__00__valueRsLineRq(x_14);
    endrule

    // No methods in this module
endmodule

interface Module188;

endinterface

module mkModule188#(function Action cache__000__setVictimRq(Struct24 _),
    function ActionValue#(Bit#(4)) getULImm_000(Struct1 _),
    function ActionValue#(Struct23) cache__000__getVictim(),
    function Action transferUpDown_000(Struct22 _),
    function Action broadcast_parentChildren000(Struct20 _),
    function Action registerDL_000(Struct19 _),
    function Action registerUL_000(Struct18 _),
    function ActionValue#(Bit#(1)) cache__000__getVictimCount(),
    function ActionValue#(Bit#(4)) getULCount_000(),
    function Action makeEnq_parentChildren000(Struct17 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__000__valueRsLineRq(Struct43 _),
    function ActionValue#(Struct13) getMSHR_000(Bit#(4) _),
    function ActionValue#(Struct42) deq_fifoL2E000(),
    function Action enq_fifoL2E000(Struct42 _),
    function ActionValue#(Struct40) cache__000__infoRsValueRq(),
    function ActionValue#(Struct3) deq_fifoI2L000(),
    function ActionValue#(Struct8) getRsReady_000(),
    function Action releaseMSHR_000(Bit#(4) _),
    function ActionValue#(Bit#(4)) cache__000__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct7) getWait_000(),
    function Action addRs_000(Struct6 _),
    function ActionValue#(Struct5) getCRqSlot_000(Struct4 _),
    function ActionValue#(Bit#(4)) findUL_000(Bit#(64) _),
    function Action enq_fifoI2L000(Struct3 _),
    function Action cache__000__infoRq(Bit#(64) _),
    function ActionValue#(Struct5) getPRqSlot_000(Struct4 _),
    function ActionValue#(Struct3) deq_fifoInput000())
    (Module188);

    rule rule_ir_prq_000;
        let x_0 <- deq_fifoInput000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_000(Struct4 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).ir_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__000__infoRq((x_2).addr);
            Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L000(x_5);
        end else begin

        end
    endrule

    rule rule_ir_prs_000;
        let x_0 <- deq_fifoInput000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- findUL_000((x_2).addr);
        let x_4 <- cache__000__infoRq((x_2).addr);
        Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : x_3});
        let x_6 <- enq_fifoI2L000(x_5);
    endrule

    rule rule_ir_crq_000;
        let x_0 <- deq_fifoInput000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getCRqSlot_000(Struct4 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__000__infoRq((x_2).addr);
            Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L000(x_5);
        end else begin

        end
    endrule

    rule rule_ir_crs_000;
        let x_0 <- deq_fifoInput000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_000(Struct6 {r_dl_midx : (x_1)[0:0], r_dl_msg :
        x_2});
    endrule

    rule rule_ir_retry_000;
        let x_0 <- getWait_000();
        when ((x_0).valid, noAction);
        Struct4 x_1 = ((x_0).data);
        Struct1 x_2 = ((x_1).r_msg);
        let x_3 <- cache__000__infoRq((x_2).addr);
        Struct3 x_4 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg : x_2,
        ir_msg_from : (x_1).r_msg_from, ir_mshr_id : (x_1).r_id});
        let x_5 <- enq_fifoI2L000(x_4);
    endrule

    rule rule_ir_invrs_000;
        let x_0 <- deq_fifoInput000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- cache__000__releaseVictim((x_2).addr);
        let x_4 <- releaseMSHR_000(x_3);
    endrule

    rule rule_ir_rsrel_000;
        let x_0 <- getRsReady_000();
        Struct1 x_1 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        let x_2 <- cache__000__infoRq((x_0).r_addr);
        Struct3 x_3 = (Struct3 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_1,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id});
        let x_4 <- enq_fifoI2L000(x_3);
    endrule

    rule rule_lr_000;
        let x_0 <- deq_fifoI2L000();
        let x_1 <- cache__000__infoRsValueRq();
        Struct42 x_2 = (Struct42 {lr_ir_pp : x_0, lr_ir : x_1});
        let x_3 <- enq_fifoL2E000(x_2);
    endrule

    rule rule_exec_000_0000000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_12).dir_st))) && ((x_11) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) :
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))}).dir_excl)))},
        value_write : (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_16}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_0010000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_010000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_000();
        let x_17 <- cache__000__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_000(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
    endrule

    rule rule_exec_000_030000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_100000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) || (((x_11) ==
        ((Bit#(3))'(3'h2))) && (((x_10) == ((Bool)'(True))) &&
        ((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) ==
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        let x_18 <- cache__000__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
    endrule

    rule rule_exec_000_110000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_000();
        let x_17 <- cache__000__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_000(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
    endrule

    rule rule_exec_000_140000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_150000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))) == ((Bit#(2))'(2'h0)))) && (((x_10) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_11))) &&
        (((x_12).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        let x_17 <- broadcast_parentChildren000(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_000_250000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren000(x_16);
    endrule

    rule rule_exec_000_26000000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_26010000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_2610000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_270000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_280000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren000(x_16);
    endrule

    rule rule_exec_000_2900000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_2910000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_2100000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_2110000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value});
        let x_19 <- cache__000__valueRsLineRq(x_18);
        Struct17 x_20 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
    endrule

    rule rule_exec_000_0400000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_0700000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_16000000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_16010000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_110000000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_110010000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_110020000;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_0000001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_12).dir_st))) && ((x_11) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) :
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))}).dir_excl)))},
        value_write : (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_16}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_0010001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_010001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_000();
        let x_17 <- cache__000__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_000(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h5))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
    endrule

    rule rule_exec_000_030001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_100001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) || (((x_11) ==
        ((Bit#(3))'(3'h2))) && (((x_10) == ((Bool)'(True))) &&
        ((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) ==
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        let x_18 <- cache__000__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
    endrule

    rule rule_exec_000_110001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_000();
        let x_17 <- cache__000__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_000(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h5))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
    endrule

    rule rule_exec_000_140001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_150001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))) == ((Bit#(2))'(2'h0)))) && (((x_10) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_11))) &&
        (((x_12).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        let x_17 <- broadcast_parentChildren000(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_000_250001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren000(x_16);
    endrule

    rule rule_exec_000_26000001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_26010001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_2610001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_270001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_280001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren000(x_16);
    endrule

    rule rule_exec_000_2900001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_2910001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_2100001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_2110001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value});
        let x_19 <- cache__000__valueRsLineRq(x_18);
        Struct17 x_20 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
    endrule

    rule rule_exec_000_0400001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_0700001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_16000001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_16010001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_110000001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_110010001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_110020001;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- addRs_000(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_000_020;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_excl)))}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_21 <- cache__000__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_000(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_24 <- makeEnq_parentChildren000(x_23);
    endrule

    rule rule_exec_000_021;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_21 <- cache__000__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_000(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_24 <- makeEnq_parentChildren000(x_23);
    endrule

    rule rule_exec_000_041;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct21 x_13 = (Struct21 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_8).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))))}, msg :
        ((x_8).m_dl_rss)[((((x_8).m_dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        (unpack(0)))))))]});
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ((x_8).m_qidx);
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : ((unpack(0)) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_st, mesi_dir_sharers : (((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        ((unpack(0)) | (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_st) ==
        ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : unpack(0), dir_sharers : ((unpack(0)) | (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0]))) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : ((unpack(0)) | (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_excl)))},
        value_write : (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (x_18).info_write, info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : (x_18).info,
        value_write : (Bool)'(True), value : ((x_13).msg).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_19).info).mesi_status,
        mesi_dir_st : ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache__000__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_000(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_14).addr, value :
        ((x_13).msg).value}});
        let x_24 <- makeEnq_parentChildren000(x_23);
    endrule

    rule rule_exec_000_05;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_12).dir_st))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_06;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_11))) && ((!
        (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_12).dir_st))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h2)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_071;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct21 x_13 = (Struct21 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_8).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))))}, msg :
        ((x_8).m_dl_rss)[((((x_8).m_dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        (unpack(0)))))))]});
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ((x_8).m_qidx);
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : (unpack(0)) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_st,
        mesi_dir_sharers : (((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        unpack(0), dir_sharers : (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : ((x_13).msg).value});
        let x_21 <- cache__000__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_000(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_14).addr, value :
        ((x_13).msg).value}});
        let x_24 <- makeEnq_parentChildren000(x_23);
    endrule

    rule rule_exec_000_12;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((((x_12).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << (({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])})[0:0])))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        let x_20 <- cache__000__valueRsLineRq(x_19);
        let x_21 <- releaseMSHR_000(x_4);
        Struct17 x_22 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
    endrule

    rule rule_exec_000_13;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])})[0:0])))) ==
        ((Bit#(2))'(2'h0)))) && (((x_12).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_15).info).mesi_status,
        mesi_dir_st : ((x_15).info).mesi_dir_st, mesi_dir_sharers :
        ((x_15).info).mesi_dir_sharers}, value_write : (x_15).value_write,
        value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        let x_18 <- transferUpDown_000(Struct22 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((x_14)[0:0])))});
        let x_19 <- broadcast_parentChildren000(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((x_14)[0:0]))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_000_161;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__000__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_000(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
    endrule

    rule rule_exec_000_170;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_171;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
    endrule

    rule rule_exec_000_190;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (x_12).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(3))'(3'h2)});
        let x_17 <- broadcast_parentChildren000(Struct20 {cs_inds :
        (x_12).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_000_191;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h2)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
    endrule

    rule rule_exec_000_192;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__000__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_000(Struct19 {r_id : x_4, r_dl_rss_from :
        (x_12).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(3))'(3'h2)});
        let x_17 <- broadcast_parentChildren000(Struct20 {cs_inds :
        (x_12).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_000_11010;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__000__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_000(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
    endrule

    rule rule_exec_000_11011;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__000__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_000(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
    endrule

    rule rule_exec_000_20;
        let x_0 <- cache__000__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_000(x_4);
        let x_6 <- cache__000__setVictimRq(Struct24 {victim_addr : x_1,
        victim_req : x_5});
        Struct13 x_7 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_9) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_10))
        && ((x_10) < ((Bit#(3))'(3'h4)))) && (((x_11).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        let x_12 <- registerUL_000(Struct18 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_14 <- makeEnq_parentChildren000(x_13);
    endrule

    rule rule_exec_000_21;
        let x_0 <- cache__000__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_000(x_4);
        let x_6 <- cache__000__setVictimRq(Struct24 {victim_addr : x_1,
        victim_req : x_5});
        Struct13 x_7 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when ((((x_11).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_9) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_10))) || (((x_9) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_10)) && ((x_10) <
        ((Bit#(3))'(3'h3)))))), noAction);
        let x_12 <- registerUL_000(Struct18 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_14 <- makeEnq_parentChildren000(x_13);
    endrule

    rule rule_exec_000_22;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h16)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when (! ((x_8).m_rsb), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__000__valueRsLineRq(x_16);
        let x_18 <- releaseMSHR_000(x_4);
    endrule

    rule rule_exec_000_23;
        let x_0 <- deq_fifoL2E000();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((((x_11) == ((Bit#(3))'(3'h1))) && (! (((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_11) == ((Bit#(3))'(3'h2))) && ((x_10)
        == ((Bool)'(False)))), noAction);
        Struct43 x_13 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_14 = (Struct43 {addr : (x_13).addr, info_write :
        (Bool)'(True), info_hit : (x_13).info_hit, info_way :
        (x_13).info_way, edir_hit : (x_13).edir_hit, edir_way :
        (x_13).edir_way, edir_slot : (x_13).edir_slot, info : Struct11
        {mesi_owned : ((x_13).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_13).info).mesi_dir_st,
        mesi_dir_sharers : ((x_13).info).mesi_dir_sharers}, value_write :
        (x_13).value_write, value : (x_13).value});
        let x_15 <- cache__000__valueRsLineRq(x_14);
    endrule

    // No methods in this module
endmodule

interface Module189;

endinterface

module mkModule189#(function Action cache__0000__setVictimRq(Struct67 _),
    function ActionValue#(Bit#(3)) getULImm_0000(Struct1 _),
    function ActionValue#(Struct66) cache__0000__getVictim(),
    function Action registerUL_0000(Struct65 _),
    function ActionValue#(Bit#(1)) cache__0000__getVictimCount(),
    function ActionValue#(Bit#(3)) getULCount_0000(),
    function Action makeEnq_parentChildren0000(Struct17 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__0000__valueRsLineRq(Struct64 _),
    function ActionValue#(Struct63) getMSHR_0000(Bit#(3) _),
    function ActionValue#(Struct62) deq_fifoL2E0000(),
    function Action enq_fifoL2E0000(Struct62 _),
    function ActionValue#(Struct60) cache__0000__infoRsValueRq(),
    function ActionValue#(Struct55) deq_fifoI2L0000(),
    function ActionValue#(Struct59) getRsReady_0000(),
    function Action releaseMSHR_0000(Bit#(3) _),
    function ActionValue#(Bit#(3)) cache__0000__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct58) getWait_0000(),
    function Action addRs_0000(Struct6 _),
    function ActionValue#(Struct57) getCRqSlot_0000(Struct56 _),
    function ActionValue#(Bit#(3)) findUL_0000(Bit#(64) _),
    function Action enq_fifoI2L0000(Struct55 _),
    function Action cache__0000__infoRq(Bit#(64) _),
    function ActionValue#(Struct57) getPRqSlot_0000(Struct56 _),
    function ActionValue#(Struct55) deq_fifoInput0000())
    (Module189);

    rule rule_ir_prq_0000;
        let x_0 <- deq_fifoInput0000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_0000(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).ir_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0000__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0000(x_5);
        end else begin

        end
    endrule

    rule rule_ir_prs_0000;
        let x_0 <- deq_fifoInput0000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- findUL_0000((x_2).addr);
        let x_4 <- cache__0000__infoRq((x_2).addr);
        Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : x_3});
        let x_6 <- enq_fifoI2L0000(x_5);
    endrule

    rule rule_ir_crq_0000;
        let x_0 <- deq_fifoInput0000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getCRqSlot_0000(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0000__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0000(x_5);
        end else begin

        end
    endrule

    rule rule_ir_crs_0000;
        let x_0 <- deq_fifoInput0000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_0000(Struct6 {r_dl_midx : (x_1)[0:0], r_dl_msg :
        x_2});
    endrule

    rule rule_ir_retry_0000;
        let x_0 <- getWait_0000();
        when ((x_0).valid, noAction);
        Struct56 x_1 = ((x_0).data);
        Struct1 x_2 = ((x_1).r_msg);
        let x_3 <- cache__0000__infoRq((x_2).addr);
        Struct55 x_4 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_2, ir_msg_from : (x_1).r_msg_from, ir_mshr_id : (x_1).r_id});
        let x_5 <- enq_fifoI2L0000(x_4);
    endrule

    rule rule_ir_invrs_0000;
        let x_0 <- deq_fifoInput0000();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- cache__0000__releaseVictim((x_2).addr);
        let x_4 <- releaseMSHR_0000(x_3);
    endrule

    rule rule_ir_rsrel_0000;
        let x_0 <- getRsReady_0000();
        Struct1 x_1 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        let x_2 <- cache__0000__infoRq((x_0).r_addr);
        Struct55 x_3 = (Struct55 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_1,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id});
        let x_4 <- enq_fifoI2L0000(x_3);
    endrule

    rule rule_lr_0000;
        let x_0 <- deq_fifoI2L0000();
        let x_1 <- cache__0000__infoRsValueRq();
        Struct62 x_2 = (Struct62 {lr_ir_pp : x_0, lr_ir : x_1});
        let x_3 <- enq_fifoL2E0000(x_2);
    endrule

    rule rule_exec_0000_00;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0000__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_15}});
        let x_17 <- makeEnq_parentChildren0000(x_16);
    endrule

    rule rule_exec_0000_01;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0000__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0000();
        let x_17 <- cache__0000__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0000(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0000(x_19);
    endrule

    rule rule_exec_0000_020;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0000__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0000(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0000(x_21);
    endrule

    rule rule_exec_0000_021;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0000__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0000(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0000(x_21);
    endrule

    rule rule_exec_0000_03;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren0000(x_18);
    endrule

    rule rule_exec_0000_100;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_11) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache__0000__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0000(x_19);
    endrule

    rule rule_exec_0000_101;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && ((x_11) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_16 <- cache__0000__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren0000(x_17);
    endrule

    rule rule_exec_0000_11;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0000__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0000();
        let x_17 <- cache__0000__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0000(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0000(x_19);
    endrule

    rule rule_exec_0000_12;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_14).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_17).info).mesi_status,
        mesi_dir_st : ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct64 x_19 = (Struct64 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        let x_20 <- cache__0000__valueRsLineRq(x_19);
        let x_21 <- releaseMSHR_0000(x_4);
        Struct17 x_22 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_23 <- makeEnq_parentChildren0000(x_22);
    endrule

    rule rule_exec_0000_130;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0000(x_18);
    endrule

    rule rule_exec_0000_131;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0000__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0000(x_18);
    endrule

    rule rule_exec_0000_20;
        let x_0 <- cache__0000__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0000(x_4);
        let x_6 <- cache__0000__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_9) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_10))
        && ((x_10) < ((Bit#(3))'(3'h4)))), noAction);
        let x_12 <- registerUL_0000(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_14 <- makeEnq_parentChildren0000(x_13);
    endrule

    rule rule_exec_0000_21;
        let x_0 <- cache__0000__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0000(x_4);
        let x_6 <- cache__0000__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_10), noAction);
        let x_12 <- registerUL_0000(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_14 <- makeEnq_parentChildren0000(x_13);
    endrule

    rule rule_exec_0000_22;
        let x_0 <- deq_fifoL2E0000();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0000(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h16)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when (! ((x_8).m_rsb), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0000__valueRsLineRq(x_16);
        let x_18 <- releaseMSHR_0000(x_4);
    endrule

    // No methods in this module
endmodule

interface Module190;

endinterface

module mkModule190#(function Action cache__0001__setVictimRq(Struct67 _),
    function ActionValue#(Bit#(3)) getULImm_0001(Struct1 _),
    function ActionValue#(Struct66) cache__0001__getVictim(),
    function Action registerUL_0001(Struct65 _),
    function ActionValue#(Bit#(1)) cache__0001__getVictimCount(),
    function ActionValue#(Bit#(3)) getULCount_0001(),
    function Action makeEnq_parentChildren0001(Struct17 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__0001__valueRsLineRq(Struct64 _),
    function ActionValue#(Struct63) getMSHR_0001(Bit#(3) _),
    function ActionValue#(Struct62) deq_fifoL2E0001(),
    function Action enq_fifoL2E0001(Struct62 _),
    function ActionValue#(Struct60) cache__0001__infoRsValueRq(),
    function ActionValue#(Struct55) deq_fifoI2L0001(),
    function ActionValue#(Struct59) getRsReady_0001(),
    function Action releaseMSHR_0001(Bit#(3) _),
    function ActionValue#(Bit#(3)) cache__0001__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct58) getWait_0001(),
    function Action addRs_0001(Struct6 _),
    function ActionValue#(Struct57) getCRqSlot_0001(Struct56 _),
    function ActionValue#(Bit#(3)) findUL_0001(Bit#(64) _),
    function Action enq_fifoI2L0001(Struct55 _),
    function Action cache__0001__infoRq(Bit#(64) _),
    function ActionValue#(Struct57) getPRqSlot_0001(Struct56 _),
    function ActionValue#(Struct55) deq_fifoInput0001())
    (Module190);

    rule rule_ir_prq_0001;
        let x_0 <- deq_fifoInput0001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_0001(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).ir_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0001__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0001(x_5);
        end else begin

        end
    endrule

    rule rule_ir_prs_0001;
        let x_0 <- deq_fifoInput0001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- findUL_0001((x_2).addr);
        let x_4 <- cache__0001__infoRq((x_2).addr);
        Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : x_3});
        let x_6 <- enq_fifoI2L0001(x_5);
    endrule

    rule rule_ir_crq_0001;
        let x_0 <- deq_fifoInput0001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getCRqSlot_0001(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0001__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0001(x_5);
        end else begin

        end
    endrule

    rule rule_ir_crs_0001;
        let x_0 <- deq_fifoInput0001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_0001(Struct6 {r_dl_midx : (x_1)[0:0], r_dl_msg :
        x_2});
    endrule

    rule rule_ir_retry_0001;
        let x_0 <- getWait_0001();
        when ((x_0).valid, noAction);
        Struct56 x_1 = ((x_0).data);
        Struct1 x_2 = ((x_1).r_msg);
        let x_3 <- cache__0001__infoRq((x_2).addr);
        Struct55 x_4 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_2, ir_msg_from : (x_1).r_msg_from, ir_mshr_id : (x_1).r_id});
        let x_5 <- enq_fifoI2L0001(x_4);
    endrule

    rule rule_ir_invrs_0001;
        let x_0 <- deq_fifoInput0001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- cache__0001__releaseVictim((x_2).addr);
        let x_4 <- releaseMSHR_0001(x_3);
    endrule

    rule rule_ir_rsrel_0001;
        let x_0 <- getRsReady_0001();
        Struct1 x_1 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        let x_2 <- cache__0001__infoRq((x_0).r_addr);
        Struct55 x_3 = (Struct55 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_1,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id});
        let x_4 <- enq_fifoI2L0001(x_3);
    endrule

    rule rule_lr_0001;
        let x_0 <- deq_fifoI2L0001();
        let x_1 <- cache__0001__infoRsValueRq();
        Struct62 x_2 = (Struct62 {lr_ir_pp : x_0, lr_ir : x_1});
        let x_3 <- enq_fifoL2E0001(x_2);
    endrule

    rule rule_exec_0001_00;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0001__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_15}});
        let x_17 <- makeEnq_parentChildren0001(x_16);
    endrule

    rule rule_exec_0001_01;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0001__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0001();
        let x_17 <- cache__0001__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0001(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0001(x_19);
    endrule

    rule rule_exec_0001_020;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0001__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0001(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0001(x_21);
    endrule

    rule rule_exec_0001_021;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0001__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0001(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0001(x_21);
    endrule

    rule rule_exec_0001_03;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren0001(x_18);
    endrule

    rule rule_exec_0001_100;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_11) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache__0001__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0001(x_19);
    endrule

    rule rule_exec_0001_101;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && ((x_11) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_16 <- cache__0001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren0001(x_17);
    endrule

    rule rule_exec_0001_11;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0001__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0001();
        let x_17 <- cache__0001__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0001(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0001(x_19);
    endrule

    rule rule_exec_0001_12;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_14).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_17).info).mesi_status,
        mesi_dir_st : ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct64 x_19 = (Struct64 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        let x_20 <- cache__0001__valueRsLineRq(x_19);
        let x_21 <- releaseMSHR_0001(x_4);
        Struct17 x_22 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_23 <- makeEnq_parentChildren0001(x_22);
    endrule

    rule rule_exec_0001_130;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0001(x_18);
    endrule

    rule rule_exec_0001_131;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0001(x_18);
    endrule

    rule rule_exec_0001_20;
        let x_0 <- cache__0001__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0001(x_4);
        let x_6 <- cache__0001__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_9) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_10))
        && ((x_10) < ((Bit#(3))'(3'h4)))), noAction);
        let x_12 <- registerUL_0001(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_14 <- makeEnq_parentChildren0001(x_13);
    endrule

    rule rule_exec_0001_21;
        let x_0 <- cache__0001__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0001(x_4);
        let x_6 <- cache__0001__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_10), noAction);
        let x_12 <- registerUL_0001(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_14 <- makeEnq_parentChildren0001(x_13);
    endrule

    rule rule_exec_0001_22;
        let x_0 <- deq_fifoL2E0001();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h16)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when (! ((x_8).m_rsb), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0001__valueRsLineRq(x_16);
        let x_18 <- releaseMSHR_0001(x_4);
    endrule

    // No methods in this module
endmodule

interface Module191;

endinterface

module mkModule191#(function Action cache__001__setVictimRq(Struct24 _),
    function ActionValue#(Bit#(4)) getULImm_001(Struct1 _),
    function ActionValue#(Struct23) cache__001__getVictim(),
    function Action transferUpDown_001(Struct22 _),
    function Action broadcast_parentChildren001(Struct20 _),
    function Action registerDL_001(Struct19 _),
    function Action registerUL_001(Struct18 _),
    function ActionValue#(Bit#(1)) cache__001__getVictimCount(),
    function ActionValue#(Bit#(4)) getULCount_001(),
    function Action makeEnq_parentChildren001(Struct17 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__001__valueRsLineRq(Struct43 _),
    function ActionValue#(Struct13) getMSHR_001(Bit#(4) _),
    function ActionValue#(Struct42) deq_fifoL2E001(),
    function Action enq_fifoL2E001(Struct42 _),
    function ActionValue#(Struct40) cache__001__infoRsValueRq(),
    function ActionValue#(Struct3) deq_fifoI2L001(),
    function ActionValue#(Struct8) getRsReady_001(),
    function Action releaseMSHR_001(Bit#(4) _),
    function ActionValue#(Bit#(4)) cache__001__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct7) getWait_001(),
    function Action addRs_001(Struct6 _),
    function ActionValue#(Struct5) getCRqSlot_001(Struct4 _),
    function ActionValue#(Bit#(4)) findUL_001(Bit#(64) _),
    function Action enq_fifoI2L001(Struct3 _),
    function Action cache__001__infoRq(Bit#(64) _),
    function ActionValue#(Struct5) getPRqSlot_001(Struct4 _),
    function ActionValue#(Struct3) deq_fifoInput001())
    (Module191);

    rule rule_ir_prq_001;
        let x_0 <- deq_fifoInput001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_001(Struct4 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).ir_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__001__infoRq((x_2).addr);
            Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L001(x_5);
        end else begin

        end
    endrule

    rule rule_ir_prs_001;
        let x_0 <- deq_fifoInput001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- findUL_001((x_2).addr);
        let x_4 <- cache__001__infoRq((x_2).addr);
        Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : x_3});
        let x_6 <- enq_fifoI2L001(x_5);
    endrule

    rule rule_ir_crq_001;
        let x_0 <- deq_fifoInput001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getCRqSlot_001(Struct4 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__001__infoRq((x_2).addr);
            Struct3 x_5 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L001(x_5);
        end else begin

        end
    endrule

    rule rule_ir_crs_001;
        let x_0 <- deq_fifoInput001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_001(Struct6 {r_dl_midx : (x_1)[0:0], r_dl_msg :
        x_2});
    endrule

    rule rule_ir_retry_001;
        let x_0 <- getWait_001();
        when ((x_0).valid, noAction);
        Struct4 x_1 = ((x_0).data);
        Struct1 x_2 = ((x_1).r_msg);
        let x_3 <- cache__001__infoRq((x_2).addr);
        Struct3 x_4 = (Struct3 {ir_is_rs_rel : (Bool)'(False), ir_msg : x_2,
        ir_msg_from : (x_1).r_msg_from, ir_mshr_id : (x_1).r_id});
        let x_5 <- enq_fifoI2L001(x_4);
    endrule

    rule rule_ir_invrs_001;
        let x_0 <- deq_fifoInput001();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- cache__001__releaseVictim((x_2).addr);
        let x_4 <- releaseMSHR_001(x_3);
    endrule

    rule rule_ir_rsrel_001;
        let x_0 <- getRsReady_001();
        Struct1 x_1 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        let x_2 <- cache__001__infoRq((x_0).r_addr);
        Struct3 x_3 = (Struct3 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_1,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id});
        let x_4 <- enq_fifoI2L001(x_3);
    endrule

    rule rule_lr_001;
        let x_0 <- deq_fifoI2L001();
        let x_1 <- cache__001__infoRsValueRq();
        Struct42 x_2 = (Struct42 {lr_ir_pp : x_0, lr_ir : x_1});
        let x_3 <- enq_fifoL2E001(x_2);
    endrule

    rule rule_exec_001_0000010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_12).dir_st))) && ((x_11) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) :
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))}).dir_excl)))},
        value_write : (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_16}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_0010010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_010010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_001();
        let x_17 <- cache__001__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_001(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
    endrule

    rule rule_exec_001_030010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_100010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) || (((x_11) ==
        ((Bit#(3))'(3'h2))) && (((x_10) == ((Bool)'(True))) &&
        ((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) ==
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        let x_18 <- cache__001__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
    endrule

    rule rule_exec_001_110010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_001();
        let x_17 <- cache__001__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_001(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
    endrule

    rule rule_exec_001_140010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_150010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))) == ((Bit#(2))'(2'h0)))) && (((x_10) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_11))) &&
        (((x_12).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h4)});
        let x_17 <- broadcast_parentChildren001(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_001_250010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren001(x_16);
    endrule

    rule rule_exec_001_26000010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_26010010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_2610010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_270010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_280010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren001(x_16);
    endrule

    rule rule_exec_001_2900010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_2910010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_2100010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h0))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h0)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_2110010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h0)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value});
        let x_19 <- cache__001__valueRsLineRq(x_18);
        Struct17 x_20 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
    endrule

    rule rule_exec_001_0400010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_0700010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_16000010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_16010010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_110000010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_110010010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_110020010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h2)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h2))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_0000011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_12).dir_st))) && ((x_11) ==
        ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) : (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) :
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))}).dir_excl)))},
        value_write : (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_16}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_0010011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_010011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_001();
        let x_17 <- cache__001__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_001(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h5))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
    endrule

    rule rule_exec_001_030011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_100011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) || (((x_11) ==
        ((Bit#(3))'(3'h2))) && (((x_10) == ((Bool)'(True))) &&
        ((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) ==
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(1))'(1'h1), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        let x_18 <- cache__001__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
    endrule

    rule rule_exec_001_110011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_11))) && (! (((Bit#(3))'(3'h2)) < ((x_12).dir_st)))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_001();
        let x_17 <- cache__001__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_001(Struct18 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h5))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
    endrule

    rule rule_exec_001_140011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_11))) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_150011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))) == ((Bit#(2))'(2'h0)))) && (((x_10) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_11))) &&
        (((x_12).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))),
        r_dl_rsb : (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h5)});
        let x_17 <- broadcast_parentChildren001(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_001_250011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren001(x_16);
    endrule

    rule rule_exec_001_26000011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_26010011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_2610011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_270011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_280011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_17 <- makeEnq_parentChildren001(x_16);
    endrule

    rule rule_exec_001_2900011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(False))) && (((((((x_12).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_2910011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(2))'(2'h1)) < ((((((x_12).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) +
        (((((((x_12).dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h1)) : ((Bit#(2))'(2'h0)))) + (unpack(0))))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl,
        dir_sharers : ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1))))}).dir_excl)))}, value_write :
        (x_14).value_write, value : (x_14).value});
        let x_16 <- cache__001__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_2100011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && (((x_11) == ((Bit#(3))'(3'h2)))
        && (((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) && (((x_12).dir_excl)
        == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1)) << ((Bit#(1))'(1'h1))))
        == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_12).dir_sharers) == (((Bit#(2))'(2'h1)) <<
        ((Bit#(1))'(1'h1)))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        ((x_14).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_14).value_write, value :
        (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_2110011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h1)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((((((x_12).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_12).dir_excl) == ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_12).dir_st) == ((Bit#(3))'(3'h3))) && (((x_12).dir_excl) ==
        ((Bit#(1))'(1'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_12).dir_sharers) | (((Bit#(2))'(2'h1))
        << ((Bit#(1))'(1'h1)))) == ((x_12).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_17).value_write, value :
        (x_17).value});
        let x_19 <- cache__001__valueRsLineRq(x_18);
        Struct17 x_20 = (Struct17 {enq_type : ((((Bit#(3))'(3'h5))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h5))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h5))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
    endrule

    rule rule_exec_001_0400011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_0700011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h6)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_16000011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_16010011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_110000011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_110010011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hf)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_110020011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h3)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hd)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- addRs_001(Struct6 {r_dl_midx : ((Bit#(3))'(3'h3))[0:0],
        r_dl_msg : x_13});
    endrule

    rule rule_exec_001_020;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_12).dir_excl, dir_sharers :
        (((x_12).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_12).dir_sharers) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) : (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0])))}).dir_excl)))}, value_write : (x_16).value_write,
        value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_21 <- cache__001__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_001(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_24 <- makeEnq_parentChildren001(x_23);
    endrule

    rule rule_exec_001_021;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_21 <- cache__001__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_001(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_24 <- makeEnq_parentChildren001(x_23);
    endrule

    rule rule_exec_001_041;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct21 x_13 = (Struct21 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_8).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))))}, msg :
        ((x_8).m_dl_rss)[((((x_8).m_dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        (unpack(0)))))))]});
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ((x_8).m_qidx);
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : ((unpack(0)) |
        (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_st, mesi_dir_sharers : (((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        ((unpack(0)) | (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_st) ==
        ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : unpack(0), dir_sharers : ((unpack(0)) | (((Bit#(2))'(2'h1)) <<
        ((x_15)[0:0]))) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : ((unpack(0)) | (((Bit#(2))'(2'h1)) << ((x_15)[0:0]))) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_excl)))},
        value_write : (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (x_18).info_write, info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : (x_18).info,
        value_write : (Bool)'(True), value : ((x_13).msg).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (Bool)'(True), info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_19).info).mesi_status,
        mesi_dir_st : ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache__001__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_001(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_14).addr, value :
        ((x_13).msg).value}});
        let x_24 <- makeEnq_parentChildren001(x_23);
    endrule

    rule rule_exec_001_05;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_12).dir_st))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_06;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_11))) && ((!
        (((x_12).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_12).dir_st))))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h3)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_071;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct21 x_13 = (Struct21 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_8).m_dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))))}, msg :
        ((x_8).m_dl_rss)[((((x_8).m_dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_8).m_dl_rss_from)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        (unpack(0)))))))]});
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ((x_8).m_qidx);
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers : (unpack(0)) |
        (((Bit#(2))'(2'h1)) << (((x_13).cidx)[0:0]))}).dir_st,
        mesi_dir_sharers : (((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        unpack(0), dir_sharers : (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15
        {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0), dir_sharers :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_sharers) : (((Bit#(2))'(2'h1)) <<
        ((Struct15 {dir_st : (Bit#(3))'(3'h2), dir_excl : unpack(0),
        dir_sharers : (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (((x_13).cidx)[0:0]))}).dir_excl)))}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        Struct43 x_20 = (Struct43 {addr : (x_19).addr, info_write :
        (x_19).info_write, info_hit : (x_19).info_hit, info_way :
        (x_19).info_way, edir_hit : (x_19).edir_hit, edir_way :
        (x_19).edir_way, edir_slot : (x_19).edir_slot, info : (x_19).info,
        value_write : (Bool)'(True), value : ((x_13).msg).value});
        let x_21 <- cache__001__valueRsLineRq(x_20);
        let x_22 <- releaseMSHR_001(x_4);
        Struct17 x_23 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_14).addr, value :
        ((x_13).msg).value}});
        let x_24 <- makeEnq_parentChildren001(x_23);
    endrule

    rule rule_exec_001_12;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((((x_12).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_12).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_12).dir_sharers) == (((Bit#(2))'(2'h1))
        << (({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])})[0:0])))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_16 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        ((x_16).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_15)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_16).value_write, value :
        (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : ((x_17).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        Struct43 x_19 = (Struct43 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_18).info).mesi_status, mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        let x_20 <- cache__001__valueRsLineRq(x_19);
        let x_21 <- releaseMSHR_001(x_4);
        Struct17 x_22 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
    endrule

    rule rule_exec_001_13;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])})[0:0])))) ==
        ((Bit#(2))'(2'h0)))) && (((x_12).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_15).info).mesi_status,
        mesi_dir_st : ((x_15).info).mesi_dir_st, mesi_dir_sharers :
        ((x_15).info).mesi_dir_sharers}, value_write : (x_15).value_write,
        value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        let x_18 <- transferUpDown_001(Struct22 {r_id : x_4, r_dl_rss_from :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((x_14)[0:0])))});
        let x_19 <- broadcast_parentChildren001(Struct20 {cs_inds :
        ((x_12).dir_sharers) & (~(((Bit#(2))'(2'h1)) << ((x_14)[0:0]))),
        cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_001_161;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_14)[0:0], dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__001__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_001(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
    endrule

    rule rule_exec_001_170;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_12).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_171;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when ((! ((x_11) < ((Bit#(3))'(3'h3)))) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
    endrule

    rule rule_exec_001_190;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (x_12).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(3))'(3'h3)});
        let x_17 <- broadcast_parentChildren001(Struct20 {cs_inds :
        (x_12).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_001_191;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && ((! (((x_12).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_12).dir_st)))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (unpack(0)) | (((Bit#(2))'(2'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_12).dir_excl)})[0:0])), r_dl_rsb :
        (Bool)'(True), r_dl_rsbTo : (Bit#(3))'(3'h3)});
        Struct17 x_17 = (Struct17 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_12).dir_excl)})[0:0], enq_msg :
        Struct1 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_13).addr, value : unpack(0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
    endrule

    rule rule_exec_001_192;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_12).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__001__valueRsLineRq(unpack(0));
        let x_16 <- registerDL_001(Struct19 {r_id : x_4, r_dl_rss_from :
        (x_12).dir_sharers, r_dl_rsb : (Bool)'(True), r_dl_rsbTo :
        (Bit#(3))'(3'h3)});
        let x_17 <- broadcast_parentChildren001(Struct20 {cs_inds :
        (x_12).dir_sharers, cs_msg : Struct1 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_13).addr, value : unpack(0)}});
    endrule

    rule rule_exec_001_11010;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__001__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_001(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
    endrule

    rule rule_exec_001_11011;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when (((x_8).m_dl_rss) == ((x_8).m_dl_rss), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = ((x_8).m_msg);
        Bit#(3) x_14 = ((x_8).m_qidx);
        Struct43 x_15 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : (Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st, mesi_dir_sharers : (((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct15 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_sharers) : (((Bit#(2))'(2'h1)) << ((Struct15 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : unpack(0), dir_sharers :
        unpack(0)}).dir_excl)))}, value_write : (x_15).value_write, value :
        (x_15).value});
        Struct43 x_17 = (Struct43 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct43 x_18 = (Struct43 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_17).info).mesi_status, mesi_dir_st : ((x_17).info).mesi_dir_st,
        mesi_dir_sharers : ((x_17).info).mesi_dir_sharers}, value_write :
        (x_17).value_write, value : (x_17).value});
        let x_19 <- cache__001__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_001(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_14)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_14)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_14)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
    endrule

    rule rule_exec_001_20;
        let x_0 <- cache__001__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_001(x_4);
        let x_6 <- cache__001__setVictimRq(Struct24 {victim_addr : x_1,
        victim_req : x_5});
        Struct13 x_7 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_9) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_10))
        && ((x_10) < ((Bit#(3))'(3'h4)))) && (((x_11).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        let x_12 <- registerUL_001(Struct18 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_14 <- makeEnq_parentChildren001(x_13);
    endrule

    rule rule_exec_001_21;
        let x_0 <- cache__001__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_001(x_4);
        let x_6 <- cache__001__setVictimRq(Struct24 {victim_addr : x_1,
        victim_req : x_5});
        Struct13 x_7 = (Struct13 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when ((((x_11).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_9) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_10))) || (((x_9) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_10)) && ((x_10) <
        ((Bit#(3))'(3'h3)))))), noAction);
        let x_12 <- registerUL_001(Struct18 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_14 <- makeEnq_parentChildren001(x_13);
    endrule

    rule rule_exec_001_22;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h16)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when (! ((x_8).m_rsb), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct43 x_14 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_15 = (Struct43 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct43 x_16 = (Struct43 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__001__valueRsLineRq(x_16);
        let x_18 <- releaseMSHR_001(x_4);
    endrule

    rule rule_exec_001_23;
        let x_0 <- deq_fifoL2E001();
        Struct3 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(4) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (x_5, noAction);
        Struct40 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_001(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((((x_11) == ((Bit#(3))'(3'h1))) && (! (((x_12).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_11) == ((Bit#(3))'(3'h2))) && ((x_10)
        == ((Bool)'(False)))), noAction);
        Struct43 x_13 = (Struct43 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct43 x_14 = (Struct43 {addr : (x_13).addr, info_write :
        (Bool)'(True), info_hit : (x_13).info_hit, info_way :
        (x_13).info_way, edir_hit : (x_13).edir_hit, edir_way :
        (x_13).edir_way, edir_slot : (x_13).edir_slot, info : Struct11
        {mesi_owned : ((x_13).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_13).info).mesi_dir_st,
        mesi_dir_sharers : ((x_13).info).mesi_dir_sharers}, value_write :
        (x_13).value_write, value : (x_13).value});
        let x_15 <- cache__001__valueRsLineRq(x_14);
    endrule

    // No methods in this module
endmodule

interface Module192;

endinterface

module mkModule192#(function Action cache__0010__setVictimRq(Struct67 _),
    function ActionValue#(Bit#(3)) getULImm_0010(Struct1 _),
    function ActionValue#(Struct66) cache__0010__getVictim(),
    function Action registerUL_0010(Struct65 _),
    function ActionValue#(Bit#(1)) cache__0010__getVictimCount(),
    function ActionValue#(Bit#(3)) getULCount_0010(),
    function Action makeEnq_parentChildren0010(Struct17 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__0010__valueRsLineRq(Struct64 _),
    function ActionValue#(Struct63) getMSHR_0010(Bit#(3) _),
    function ActionValue#(Struct62) deq_fifoL2E0010(),
    function Action enq_fifoL2E0010(Struct62 _),
    function ActionValue#(Struct60) cache__0010__infoRsValueRq(),
    function ActionValue#(Struct55) deq_fifoI2L0010(),
    function ActionValue#(Struct59) getRsReady_0010(),
    function Action releaseMSHR_0010(Bit#(3) _),
    function ActionValue#(Bit#(3)) cache__0010__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct58) getWait_0010(),
    function Action addRs_0010(Struct6 _),
    function ActionValue#(Struct57) getCRqSlot_0010(Struct56 _),
    function ActionValue#(Bit#(3)) findUL_0010(Bit#(64) _),
    function Action enq_fifoI2L0010(Struct55 _),
    function Action cache__0010__infoRq(Bit#(64) _),
    function ActionValue#(Struct57) getPRqSlot_0010(Struct56 _),
    function ActionValue#(Struct55) deq_fifoInput0010())
    (Module192);

    rule rule_ir_prq_0010;
        let x_0 <- deq_fifoInput0010();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_0010(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).ir_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0010__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0010(x_5);
        end else begin

        end
    endrule

    rule rule_ir_prs_0010;
        let x_0 <- deq_fifoInput0010();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- findUL_0010((x_2).addr);
        let x_4 <- cache__0010__infoRq((x_2).addr);
        Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : x_3});
        let x_6 <- enq_fifoI2L0010(x_5);
    endrule

    rule rule_ir_crq_0010;
        let x_0 <- deq_fifoInput0010();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getCRqSlot_0010(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0010__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0010(x_5);
        end else begin

        end
    endrule

    rule rule_ir_crs_0010;
        let x_0 <- deq_fifoInput0010();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_0010(Struct6 {r_dl_midx : (x_1)[0:0], r_dl_msg :
        x_2});
    endrule

    rule rule_ir_retry_0010;
        let x_0 <- getWait_0010();
        when ((x_0).valid, noAction);
        Struct56 x_1 = ((x_0).data);
        Struct1 x_2 = ((x_1).r_msg);
        let x_3 <- cache__0010__infoRq((x_2).addr);
        Struct55 x_4 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_2, ir_msg_from : (x_1).r_msg_from, ir_mshr_id : (x_1).r_id});
        let x_5 <- enq_fifoI2L0010(x_4);
    endrule

    rule rule_ir_invrs_0010;
        let x_0 <- deq_fifoInput0010();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- cache__0010__releaseVictim((x_2).addr);
        let x_4 <- releaseMSHR_0010(x_3);
    endrule

    rule rule_ir_rsrel_0010;
        let x_0 <- getRsReady_0010();
        Struct1 x_1 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        let x_2 <- cache__0010__infoRq((x_0).r_addr);
        Struct55 x_3 = (Struct55 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_1,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id});
        let x_4 <- enq_fifoI2L0010(x_3);
    endrule

    rule rule_lr_0010;
        let x_0 <- deq_fifoI2L0010();
        let x_1 <- cache__0010__infoRsValueRq();
        Struct62 x_2 = (Struct62 {lr_ir_pp : x_0, lr_ir : x_1});
        let x_3 <- enq_fifoL2E0010(x_2);
    endrule

    rule rule_exec_0010_00;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0010__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_15}});
        let x_17 <- makeEnq_parentChildren0010(x_16);
    endrule

    rule rule_exec_0010_01;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0010__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0010();
        let x_17 <- cache__0010__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0010(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0010(x_19);
    endrule

    rule rule_exec_0010_020;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0010__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0010(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0010(x_21);
    endrule

    rule rule_exec_0010_021;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0010__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0010(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0010(x_21);
    endrule

    rule rule_exec_0010_03;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0010__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren0010(x_18);
    endrule

    rule rule_exec_0010_100;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_11) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache__0010__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0010(x_19);
    endrule

    rule rule_exec_0010_101;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && ((x_11) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_16 <- cache__0010__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren0010(x_17);
    endrule

    rule rule_exec_0010_11;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0010__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0010();
        let x_17 <- cache__0010__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0010(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0010(x_19);
    endrule

    rule rule_exec_0010_12;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_14).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_17).info).mesi_status,
        mesi_dir_st : ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct64 x_19 = (Struct64 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        let x_20 <- cache__0010__valueRsLineRq(x_19);
        let x_21 <- releaseMSHR_0010(x_4);
        Struct17 x_22 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_23 <- makeEnq_parentChildren0010(x_22);
    endrule

    rule rule_exec_0010_130;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0010__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0010(x_18);
    endrule

    rule rule_exec_0010_131;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h4)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0010__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h2))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h2))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h2))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0010(x_18);
    endrule

    rule rule_exec_0010_20;
        let x_0 <- cache__0010__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0010(x_4);
        let x_6 <- cache__0010__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_9) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_10))
        && ((x_10) < ((Bit#(3))'(3'h4)))), noAction);
        let x_12 <- registerUL_0010(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_14 <- makeEnq_parentChildren0010(x_13);
    endrule

    rule rule_exec_0010_21;
        let x_0 <- cache__0010__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0010(x_4);
        let x_6 <- cache__0010__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_10), noAction);
        let x_12 <- registerUL_0010(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h0))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h0))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h0))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_14 <- makeEnq_parentChildren0010(x_13);
    endrule

    rule rule_exec_0010_22;
        let x_0 <- deq_fifoL2E0010();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0010(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h0))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h16)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when (! ((x_8).m_rsb), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0010__valueRsLineRq(x_16);
        let x_18 <- releaseMSHR_0010(x_4);
    endrule

    // No methods in this module
endmodule

interface Module193;

endinterface

module mkModule193#(function Action cache__0011__setVictimRq(Struct67 _),
    function ActionValue#(Bit#(3)) getULImm_0011(Struct1 _),
    function ActionValue#(Struct66) cache__0011__getVictim(),
    function Action registerUL_0011(Struct65 _),
    function ActionValue#(Bit#(1)) cache__0011__getVictimCount(),
    function ActionValue#(Bit#(3)) getULCount_0011(),
    function Action makeEnq_parentChildren0011(Struct17 _),
    function ActionValue#(Vector#(4, Bit#(64))) cache__0011__valueRsLineRq(Struct64 _),
    function ActionValue#(Struct63) getMSHR_0011(Bit#(3) _),
    function ActionValue#(Struct62) deq_fifoL2E0011(),
    function Action enq_fifoL2E0011(Struct62 _),
    function ActionValue#(Struct60) cache__0011__infoRsValueRq(),
    function ActionValue#(Struct55) deq_fifoI2L0011(),
    function ActionValue#(Struct59) getRsReady_0011(),
    function Action releaseMSHR_0011(Bit#(3) _),
    function ActionValue#(Bit#(3)) cache__0011__releaseVictim(Bit#(64) _),
    function ActionValue#(Struct58) getWait_0011(),
    function Action addRs_0011(Struct6 _),
    function ActionValue#(Struct57) getCRqSlot_0011(Struct56 _),
    function ActionValue#(Bit#(3)) findUL_0011(Bit#(64) _),
    function Action enq_fifoI2L0011(Struct55 _),
    function Action cache__0011__infoRq(Bit#(64) _),
    function ActionValue#(Struct57) getPRqSlot_0011(Struct56 _),
    function ActionValue#(Struct55) deq_fifoInput0011())
    (Module193);

    rule rule_ir_prq_0011;
        let x_0 <- deq_fifoInput0011();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getPRqSlot_0011(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : (x_0).ir_msg_from});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0011__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0011(x_5);
        end else begin

        end
    endrule

    rule rule_ir_prs_0011;
        let x_0 <- deq_fifoInput0011();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (! (((x_2).id) == ((Bit#(6))'(6'h16)))),
        noAction);
        let x_3 <- findUL_0011((x_2).addr);
        let x_4 <- cache__0011__infoRq((x_2).addr);
        Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : x_3});
        let x_6 <- enq_fifoI2L0011(x_5);
    endrule

    rule rule_ir_crq_0011;
        let x_0 <- deq_fifoInput0011();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h0)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (! ((x_2).type_), noAction);
        let x_3 <- getCRqSlot_0011(Struct56 {r_id : unpack(0), r_msg : x_2,
        r_msg_from : x_1});
        when ((x_3).s_has_slot,
        noAction);
        if (! ((x_3).s_conflict)) begin
            let x_4 <- cache__0011__infoRq((x_2).addr);
            Struct55 x_5 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
            (x_0).ir_msg, ir_msg_from : x_1, ir_mshr_id : (x_3).s_id});
            let x_6 <- enq_fifoI2L0011(x_5);
        end else begin

        end
    endrule

    rule rule_ir_crs_0011;
        let x_0 <- deq_fifoInput0011();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when (((x_1)[2:1]) == ((Bit#(2))'(2'h1)), noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when ((x_2).type_, noAction);
        let x_3 <- addRs_0011(Struct6 {r_dl_midx : (x_1)[0:0], r_dl_msg :
        x_2});
    endrule

    rule rule_ir_retry_0011;
        let x_0 <- getWait_0011();
        when ((x_0).valid, noAction);
        Struct56 x_1 = ((x_0).data);
        Struct1 x_2 = ((x_1).r_msg);
        let x_3 <- cache__0011__infoRq((x_2).addr);
        Struct55 x_4 = (Struct55 {ir_is_rs_rel : (Bool)'(False), ir_msg :
        x_2, ir_msg_from : (x_1).r_msg_from, ir_mshr_id : (x_1).r_id});
        let x_5 <- enq_fifoI2L0011(x_4);
    endrule

    rule rule_ir_invrs_0011;
        let x_0 <- deq_fifoInput0011();
        Bit#(3) x_1 = ((x_0).ir_msg_from);
        when ((x_1) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        Struct1 x_2 = ((x_0).ir_msg);
        when (((x_2).type_) && (((x_2).id) == ((Bit#(6))'(6'h16))),
        noAction);
        let x_3 <- cache__0011__releaseVictim((x_2).addr);
        let x_4 <- releaseMSHR_0011(x_3);
    endrule

    rule rule_ir_rsrel_0011;
        let x_0 <- getRsReady_0011();
        Struct1 x_1 = (Struct1 {id : unpack(0), type_ : unpack(0), addr :
        (x_0).r_addr, value : unpack(0)});
        let x_2 <- cache__0011__infoRq((x_0).r_addr);
        Struct55 x_3 = (Struct55 {ir_is_rs_rel : (Bool)'(True), ir_msg : x_1,
        ir_msg_from : unpack(0), ir_mshr_id : (x_0).r_id});
        let x_4 <- enq_fifoI2L0011(x_3);
    endrule

    rule rule_lr_0011;
        let x_0 <- deq_fifoI2L0011();
        let x_1 <- cache__0011__infoRsValueRq();
        Struct62 x_2 = (Struct62 {lr_ir_pp : x_0, lr_ir : x_1});
        let x_3 <- enq_fifoL2E0011(x_2);
    endrule

    rule rule_exec_0011_00;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0011__valueRsLineRq(unpack(0));
        Struct17 x_16 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_15}});
        let x_17 <- makeEnq_parentChildren0011(x_16);
    endrule

    rule rule_exec_0011_01;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0011__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0011();
        let x_17 <- cache__0011__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0011(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0011(x_19);
    endrule

    rule rule_exec_0011_020;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h3)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0011__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0011(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0011(x_21);
    endrule

    rule rule_exec_0011_021;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h4)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : ((x_16).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h3), mesi_dir_st : ((x_16).info).mesi_dir_st,
        mesi_dir_sharers : ((x_16).info).mesi_dir_sharers}, value_write :
        (x_16).value_write, value : (x_16).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (x_17).info_write, info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : (x_17).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_19 <- cache__0011__valueRsLineRq(x_18);
        let x_20 <- releaseMSHR_0011(x_4);
        Struct17 x_21 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_13).addr, value :
        (x_13).value}});
        let x_22 <- makeEnq_parentChildren0011(x_21);
    endrule

    rule rule_exec_0011_03;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h2))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h2), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0011__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_13).addr, value :
        x_17}});
        let x_19 <- makeEnq_parentChildren0011(x_18);
    endrule

    rule rule_exec_0011_100;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when ((x_11) == ((Bit#(3))'(3'h3)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : ((x_15).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (Bool)'(True), info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_16).info).mesi_status,
        mesi_dir_st : ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache__0011__valueRsLineRq(x_17);
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0011(x_19);
    endrule

    rule rule_exec_0011_101;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (((x_10) == ((Bool)'(True))) && ((x_11) == ((Bit#(3))'(3'h4))),
        noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (x_14).info_write, info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : (x_14).info,
        value_write : (Bool)'(True), value : (x_13).value});
        let x_16 <- cache__0011__valueRsLineRq(x_15);
        Struct17 x_17 = (Struct17 {enq_type : ((((Bit#(3))'(3'h4))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h4))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h4))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_18 <- makeEnq_parentChildren0011(x_17);
    endrule

    rule rule_exec_0011_11;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_3).type_), noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_11)), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        let x_15 <- cache__0011__valueRsLineRq(unpack(0));
        let x_16 <- getULCount_0011();
        let x_17 <- cache__0011__getVictimCount();
        when ((x_16) < (zeroExtend(-(x_17))), noAction);
        let x_18 <- registerUL_0011(Struct65 {r_id : x_4, r_ul_rsb :
        (Bool)'(True), r_ul_rsbTo : ((Bit#(3))'(3'h4))[0:0]});
        Struct17 x_19 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_13).addr, value :
        unpack(0)}});
        let x_20 <- makeEnq_parentChildren0011(x_19);
    endrule

    rule rule_exec_0011_12;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hb)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((((x_8).m_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_8).m_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when ((x_8).m_rsb, noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct1 x_14 = ((x_8).m_msg);
        Bit#(3) x_15 = ({((Bit#(2))'(2'h2)),(((x_8).m_qidx)[0:0])});
        Struct64 x_16 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_17 = (Struct64 {addr : (x_16).addr, info_write :
        (x_16).info_write, info_hit : (x_16).info_hit, info_way :
        (x_16).info_way, edir_hit : (x_16).edir_hit, edir_way :
        (x_16).edir_way, edir_slot : (x_16).edir_slot, info : (x_16).info,
        value_write : (Bool)'(True), value : (x_14).value});
        Struct64 x_18 = (Struct64 {addr : (x_17).addr, info_write :
        (Bool)'(True), info_hit : (x_17).info_hit, info_way :
        (x_17).info_way, edir_hit : (x_17).edir_hit, edir_way :
        (x_17).edir_way, edir_slot : (x_17).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(True), mesi_status : ((x_17).info).mesi_status,
        mesi_dir_st : ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct64 x_19 = (Struct64 {addr : (x_18).addr, info_write :
        (Bool)'(True), info_hit : (x_18).info_hit, info_way :
        (x_18).info_way, edir_hit : (x_18).edir_hit, edir_way :
        (x_18).edir_way, edir_slot : (x_18).edir_slot, info : Struct11
        {mesi_owned : ((x_18).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h4), mesi_dir_st : ((x_18).info).mesi_dir_st,
        mesi_dir_sharers : ((x_18).info).mesi_dir_sharers}, value_write :
        (x_18).value_write, value : (x_18).value});
        let x_20 <- cache__0011__valueRsLineRq(x_19);
        let x_21 <- releaseMSHR_0011(x_4);
        Struct17 x_22 = (Struct17 {enq_type : (((x_15)[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_15)[2:1]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_15)[0:0], enq_msg : Struct1 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_13).addr, value : unpack(0)}});
        let x_23 <- makeEnq_parentChildren0011(x_22);
    endrule

    rule rule_exec_0011_130;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_3).type_), noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0011__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0011(x_18);
    endrule

    rule rule_exec_0011_131;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ((Bit#(3))'(3'h5)), noAction);
        when (((x_3).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_3).type_), noAction);
        when (! ((x_11) < ((Bit#(3))'(3'h3))), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h1), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0011__valueRsLineRq(x_16);
        Struct17 x_18 = (Struct17 {enq_type : ((((Bit#(3))'(3'h3))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h3))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h3))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_13).addr, value :
        unpack(0)}});
        let x_19 <- makeEnq_parentChildren0011(x_18);
    endrule

    rule rule_exec_0011_20;
        let x_0 <- cache__0011__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0011(x_4);
        let x_6 <- cache__0011__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((x_9) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_10))
        && ((x_10) < ((Bit#(3))'(3'h4)))), noAction);
        let x_12 <- registerUL_0011(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_4).addr, value :
        unpack(0)}});
        let x_14 <- makeEnq_parentChildren0011(x_13);
    endrule

    rule rule_exec_0011_21;
        let x_0 <- cache__0011__getVictim();
        Bit#(64) x_1 = ((x_0).victim_addr);
        Struct11 x_2 = ((x_0).victim_info);
        Vector#(4, Bit#(64)) x_3 = ((x_0).victim_value);
        Struct1 x_4 = (Struct1 {id : unpack(0), type_ : (Bool)'(False), addr
        : x_1, value : unpack(0)});
        let x_5 <- getULImm_0011(x_4);
        let x_6 <- cache__0011__setVictimRq(Struct67 {victim_addr : x_1,
        victim_req : x_5});
        Struct63 x_7 = (Struct63 {m_status : (Bit#(2))'(2'h3), m_next :
        unpack(0), m_is_ul : (Bool)'(True), m_msg : x_4, m_qidx : unpack(0),
        m_rsb : (Bool)'(False), m_dl_rss_from : unpack(0), m_dl_rss_recv :
        unpack(0), m_dl_rss : unpack(0)});
        Vector#(4, Bit#(64)) x_8 = (unpack(0));
        Bool x_9 = ((x_2).mesi_owned);
        Bit#(3) x_10 = ((x_2).mesi_status);
        Struct15 x_11 = (Struct15 {dir_st : (x_2).mesi_dir_st, dir_excl :
        ((((x_2).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_2).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_2).mesi_dir_sharers});
        when (! ((x_4).type_), noAction);
        when (((Bit#(3))'(3'h0)) < (x_10), noAction);
        let x_12 <- registerUL_0011(Struct65 {r_id : x_5, r_ul_rsb :
        (Bool)'(False), r_ul_rsbTo : unpack(0)});
        Struct17 x_13 = (Struct17 {enq_type : ((((Bit#(3))'(3'h1))[2:1]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(3))'(3'h1))[2:1])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(3))'(3'h1))[0:0], enq_msg : Struct1 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_4).addr, value :
        x_3}});
        let x_14 <- makeEnq_parentChildren0011(x_13);
    endrule

    rule rule_exec_0011_22;
        let x_0 <- deq_fifoL2E0011();
        Struct55 x_1 = ((x_0).lr_ir_pp);
        Bit#(3) x_2 = ((x_1).ir_msg_from);
        Struct1 x_3 = ((x_1).ir_msg);
        Bit#(3) x_4 = ((x_1).ir_mshr_id);
        Bool x_5 = ((x_1).ir_is_rs_rel);
        when (! (x_5), noAction);
        Struct60 x_6 = ((x_0).lr_ir);
        Struct11 x_7 = ((x_6).info);
        let x_8 <- getMSHR_0011(x_4);
        Vector#(4, Bit#(64)) x_9 = (unpack(0));
        Bool x_10 = ((x_7).mesi_owned);
        Bit#(3) x_11 = ((x_7).mesi_status);
        Struct15 x_12 = (Struct15 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) +
        ((((((x_7).mesi_dir_sharers)[1:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(1))'(1'h0)) : (((Bit#(1))'(1'h1)) + (unpack(0))))))),
        dir_sharers : (x_7).mesi_dir_sharers});
        when ((x_2) == ({((Bit#(2))'(2'h2)),((Bit#(1))'(1'h1))}),
        noAction);
        when (((x_3).id) == ((Bit#(6))'(6'h16)), noAction);
        when (((x_8).m_status) == ((Bit#(2))'(2'h3)), noAction);
        when (! ((x_8).m_rsb), noAction);
        when ((x_3).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct1 x_13 = (x_3);
        Struct64 x_14 = (Struct64 {addr : (x_3).addr, info_write :
        (Bool)'(False), info_hit : (x_6).info_hit, info_way : (x_6).info_way,
        edir_hit : (x_6).edir_hit, edir_way : (x_6).edir_way, edir_slot :
        (x_6).edir_slot, info : (x_6).info, value_write : (Bool)'(False),
        value : unpack(0)});
        Struct64 x_15 = (Struct64 {addr : (x_14).addr, info_write :
        (Bool)'(True), info_hit : (x_14).info_hit, info_way :
        (x_14).info_way, edir_hit : (x_14).edir_hit, edir_way :
        (x_14).edir_way, edir_slot : (x_14).edir_slot, info : Struct11
        {mesi_owned : ((x_14).info).mesi_owned, mesi_status :
        (Bit#(3))'(3'h0), mesi_dir_st : ((x_14).info).mesi_dir_st,
        mesi_dir_sharers : ((x_14).info).mesi_dir_sharers}, value_write :
        (x_14).value_write, value : (x_14).value});
        Struct64 x_16 = (Struct64 {addr : (x_15).addr, info_write :
        (Bool)'(True), info_hit : (x_15).info_hit, info_way :
        (x_15).info_way, edir_hit : (x_15).edir_hit, edir_way :
        (x_15).edir_way, edir_slot : (x_15).edir_slot, info : Struct11
        {mesi_owned : (Bool)'(False), mesi_status :
        ((x_15).info).mesi_status, mesi_dir_st : ((x_15).info).mesi_dir_st,
        mesi_dir_sharers : ((x_15).info).mesi_dir_sharers}, value_write :
        (x_15).value_write, value : (x_15).value});
        let x_17 <- cache__0011__valueRsLineRq(x_16);
        let x_18 <- releaseMSHR_0011(x_4);
    endrule

    // No methods in this module
endmodule

// The CC interface is defined in the header part (thus in Header.bsv)

module mkCC#(function ActionValue#(Struct1) deq_fifo002(),
function Action enq_fifo001(Struct1 _),
function Action enq_fifo000(Struct1 _)) (CC);
    Module1 m1 <- mkModule1 ();
    Module2 m2 <- mkModule2 ();
    Module3 m3 <- mkModule3 ();
    Module4 m4 <- mkModule4 ();
    Module5 m5 <- mkModule5 ();
    Module6 m6 <- mkModule6 ();
    Module7 m7 <- mkModule7 ();
    Module8 m8 <- mkModule8 ();
    Module9 m9 <- mkModule9 ();
    Module10 m10 <- mkModule10 ();
    Module11 m11 <- mkModule11 ();
    Module12 m12 <- mkModule12 ();
    Module13 m13 <- mkModule13 ();
    Module14 m14 <- mkModule14 ();
    Module15 m15 <- mkModule15 ();
    Module16 m16 <- mkModule16 ();
    Module17 m17 <- mkModule17 ();
    Module18 m18 <- mkModule18 ();
    Module19 m19 <- mkModule19 ();
    Module20 m20 <- mkModule20 ();
    Module21 m21 <- mkModule21 ();
    Module22 m22 <- mkModule22 ();
    Module23 m23 <- mkModule23 ();
    Module24 m24 <- mkModule24 ();
    Module25 m25 <- mkModule25 ();
    Module26 m26 <- mkModule26 ();
    Module27 m27 <- mkModule27 ();
    Module28 m28 <- mkModule28 ();
    Module29 m29 <- mkModule29 ();
    Module30 m30 <- mkModule30 ();
    Module31 m31 <- mkModule31 ();
    Module32 m32 <- mkModule32 ();
    Module33 m33 <- mkModule33 ();
    Module34 m34 <- mkModule34 ();
    Module35 m35 <- mkModule35 ();
    Module36 m36 <- mkModule36 ();
    Module37 m37 <- mkModule37 ();
    Module38 m38 <- mkModule38 ();
    Module39 m39 <- mkModule39 ();
    Module40 m40 <- mkModule40 ();
    Module41 m41 <- mkModule41 ();
    Module42 m42 <- mkModule42 ();
    Module43 m43 <- mkModule43 ();
    Module44 m44 <- mkModule44 ();
    Module45 m45 <- mkModule45 ();
    Module46 m46 <- mkModule46 ();
    Module47 m47 <- mkModule47 ();
    Module48 m48 <- mkModule48 ();
    Module49 m49 <- mkModule49 ();
    Module50 m50 <- mkModule50 ();
    Module51 m51 <- mkModule51 ();
    Module52 m52 <- mkModule52 ();
    Module53 m53 <- mkModule53 ();
    Module54 m54 <- mkModule54 ();
    Module55 m55 <- mkModule55 ();
    Module56 m56 <- mkModule56 ();
    Module57 m57 <- mkModule57 ();
    Module58 m58 <- mkModule58 ();
    Module59 m59 <- mkModule59 ();
    Module60 m60 <- mkModule60 ();
    Module61 m61 <- mkModule61 ();
    Module62 m62 <- mkModule62 ();
    Module63 m63 <- mkModule63 ();
    Module64 m64 <- mkModule64 ();
    Module65 m65 <- mkModule65 ();
    Module66 m66 <- mkModule66 ();
    Module67 m67 <- mkModule67 ();
    Module68 m68 <- mkModule68 ();
    Module69 m69 <- mkModule69 ();
    Module70 m70 <- mkModule70 ();
    Module71 m71 <- mkModule71 ();
    Module72 m72 <- mkModule72 ();
    Module73 m73 <- mkModule73 ();
    Module74 m74 <- mkModule74 ();
    Module75 m75 <- mkModule75 ();
    Module76 m76 <- mkModule76 ();
    Module77 m77 <- mkModule77 ();
    Module78 m78 <- mkModule78 ();
    Module79 m79 <- mkModule79 ();
    Module80 m80 <- mkModule80 ();
    Module81 m81 <- mkModule81 ();
    Module82 m82 <- mkModule82 ();
    Module83 m83 <- mkModule83 ();
    Module84 m84 <- mkModule84 ();
    Module85 m85 <- mkModule85 ();
    Module86 m86 <- mkModule86 ();
    Module87 m87 <- mkModule87 ();
    Module88 m88 <- mkModule88 ();
    Module89 m89 <- mkModule89 ();
    Module90 m90 <- mkModule90 ();
    Module91 m91 <- mkModule91 ();
    Module92 m92 <- mkModule92 ();
    Module93 m93 <- mkModule93 ();
    Module94 m94 <- mkModule94 ();
    Module95 m95 <- mkModule95 ();
    Module96 m96 <- mkModule96 ();
    Module97 m97 <- mkModule97 ();
    Module98 m98 <- mkModule98 ();
    Module99 m99 <- mkModule99 ();
    Module100 m100 <- mkModule100 ();
    Module101 m101 <- mkModule101 ();
    Module102 m102 <- mkModule102 ();
    Module103 m103 <- mkModule103 ();
    Module104 m104 <- mkModule104 ();
    Module105 m105 <- mkModule105 ();
    Module106 m106 <- mkModule106 ();
    Module107 m107 <- mkModule107 ();
    Module108 m108 <- mkModule108 ();
    Module109 m109 <- mkModule109 ();
    Module110 m110 <- mkModule110 ();
    Module111 m111 <- mkModule111 ();
    Module112 m112 <- mkModule112 ();
    Module113 m113 <- mkModule113 ();
    Module114 m114 <- mkModule114 ();
    Module115 m115 <- mkModule115 ();
    Module116 m116 <- mkModule116 ();
    Module117 m117 <- mkModule117 ();
    Module118 m118 <- mkModule118 ();
    Module119 m119 <- mkModule119 ();
    Module120 m120 <- mkModule120 ();
    Module121 m121 <- mkModule121 ();
    Module122 m122 <- mkModule122 ();
    Module123 m123 <- mkModule123 ();
    Module124 m124 <- mkModule124 ();
    Module125 m125 <- mkModule125 ();
    Module126 m126 <- mkModule126 ();
    Module127 m127 <- mkModule127 ();
    Module128 m128 <- mkModule128 ();
    Module129 m129 <- mkModule129 ();
    Module130 m130 <- mkModule130 ();
    Module131 m131 <- mkModule131 ();
    Module132 m132 <- mkModule132 ();
    Module133 m133 <- mkModule133 ();
    Module134 m134 <- mkModule134 ();
    Module135 m135 <- mkModule135 ();
    Module136 m136 <- mkModule136 ();
    Module137 m137 <- mkModule137 ();
    Module138 m138 <- mkModule138 ();
    Module139 m139 <- mkModule139 ();
    Module140 m140 <- mkModule140 ();
    Module141 m141 <- mkModule141 ();
    Module142 m142 <- mkModule142 ();
    Module143 m143 <- mkModule143 ();
    Module144 m144 <- mkModule144 ();
    Module145 m145 <- mkModule145 ();
    Module146 m146 <- mkModule146 ();
    Module147 m147 <- mkModule147 ();
    Module148 m148 <- mkModule148 ();
    Module149 m149 <- mkModule149 ();
    Module150 m150 <- mkModule150 ();
    Module151 m151 <- mkModule151 ();
    Module152 m152 <- mkModule152 ();
    Module153 m153 <- mkModule153 (m99.deq_fifo0010, m1.enq_fifoCRqInput00,
    m40.deq_fifo0000);
    Module154 m154 <- mkModule154 (m99.deq_fifo0010, m2.enq_fifoCRsInput00,
    m40.deq_fifo0000);
    Module155 m155 <- mkModule155 (m2.deq_fifoCRsInput00,
    m1.deq_fifoCRqInput00, m3.enq_fifoInput00, deq_fifo002);
    Module156 m156 <- mkModule156 (m42.enq_fifo0002, m101.enq_fifo0012,
    enq_fifo001, enq_fifo000);
    Module157 m157 <- mkModule157 (m33.wrReq_repRam__00,
    m33.rdResp_repRam__00, m33.rdReq_repRam__00);
    Module158 m158 <- mkModule158 (m80.deq_fifo00010,
    m35.enq_fifoCRqInput000, m63.deq_fifo00000);
    Module159 m159 <- mkModule159 (m80.deq_fifo00010,
    m36.enq_fifoCRsInput000, m63.deq_fifo00000);
    Module160 m160 <- mkModule160 (m36.deq_fifoCRsInput000,
    m35.deq_fifoCRqInput000, m37.enq_fifoInput000, m42.deq_fifo0002);

    Module161 m161 <- mkModule161 (m65.enq_fifo00002, m82.enq_fifo00012,
    m41.enq_fifo0001, m40.enq_fifo0000);
    Module162 m162 <- mkModule162 (m58.wrReq_repRam__000,
    m58.rdResp_repRam__000, m58.rdReq_repRam__000);
    Module163 m163 <- mkModule163 (m66.deq_fifo000000, m60.enq_fifoInput0000,
    m65.deq_fifo00002);
    Module164 m164 <- mkModule164 (m67.enq_fifo000002, m64.enq_fifo00001,
    m63.enq_fifo00000);
    Module165 m165 <- mkModule165 (m75.wrReq_repRam__0000,
    m75.rdResp_repRam__0000, m75.rdReq_repRam__0000);
    Module166 m166 <- mkModule166 (m83.deq_fifo000100, m77.enq_fifoInput0001,
    m82.deq_fifo00012);
    Module167 m167 <- mkModule167 (m84.enq_fifo000102, m81.enq_fifo00011,
    m80.enq_fifo00010);
    Module168 m168 <- mkModule168 (m92.wrReq_repRam__0001,
    m92.rdResp_repRam__0001, m92.rdReq_repRam__0001);
    Module169 m169 <- mkModule169 (m139.deq_fifo00110,
    m94.enq_fifoCRqInput001, m122.deq_fifo00100);
    Module170 m170 <- mkModule170 (m139.deq_fifo00110,
    m95.enq_fifoCRsInput001, m122.deq_fifo00100);
    Module171 m171 <- mkModule171 (m95.deq_fifoCRsInput001,
    m94.deq_fifoCRqInput001, m96.enq_fifoInput001, m101.deq_fifo0012);

    Module172 m172 <- mkModule172 (m124.enq_fifo00102, m141.enq_fifo00112,
    m100.enq_fifo0011, m99.enq_fifo0010);
    Module173 m173 <- mkModule173 (m117.wrReq_repRam__001,
    m117.rdResp_repRam__001, m117.rdReq_repRam__001);
    Module174 m174 <- mkModule174 (m125.deq_fifo001000,
    m119.enq_fifoInput0010, m124.deq_fifo00102);
    Module175 m175 <- mkModule175 (m126.enq_fifo001002, m123.enq_fifo00101,
    m122.enq_fifo00100);
    Module176 m176 <- mkModule176 (m134.wrReq_repRam__0010,
    m134.rdResp_repRam__0010, m134.rdReq_repRam__0010);
    Module177 m177 <- mkModule177 (m142.deq_fifo001100,
    m136.enq_fifoInput0011, m141.deq_fifo00112);
    Module178 m178 <- mkModule178 (m143.enq_fifo001102, m140.enq_fifo00111,
    m139.enq_fifo00110);
    Module179 m179 <- mkModule179 (m151.wrReq_repRam__0011,
    m151.rdResp_repRam__0011, m151.rdReq_repRam__0011);
    Module180 m180 <- mkModule180 (m24.wrReq_edirRam__00__7,
    m25.wrReq_edirRam__00__6, m26.wrReq_edirRam__00__5,
    m27.wrReq_edirRam__00__4, m28.wrReq_edirRam__00__3,
    m29.wrReq_edirRam__00__2, m30.wrReq_edirRam__00__1,
    m31.wrReq_edirRam__00__0, m32.wrReq_dataRam__00, m157.repAccess__00,
    m8.wrReq_infoRam__00__15, m9.wrReq_infoRam__00__14,
    m10.wrReq_infoRam__00__13, m11.wrReq_infoRam__00__12,
    m12.wrReq_infoRam__00__11, m13.wrReq_infoRam__00__10,
    m14.wrReq_infoRam__00__9, m15.wrReq_infoRam__00__8,
    m16.wrReq_infoRam__00__7, m17.wrReq_infoRam__00__6,
    m18.wrReq_infoRam__00__5, m19.wrReq_infoRam__00__4,
    m20.wrReq_infoRam__00__3, m21.wrReq_infoRam__00__2,
    m22.wrReq_infoRam__00__1, m23.wrReq_infoRam__00__0,
    m32.rdResp_dataRam__00, m7.deq_cp_2__00, m32.rdReq_dataRam__00,
    m157.repGetRs__00, m24.rdResp_edirRam__00__7, m25.rdResp_edirRam__00__6,
    m26.rdResp_edirRam__00__5, m27.rdResp_edirRam__00__4,
    m28.rdResp_edirRam__00__3, m29.rdResp_edirRam__00__2,
    m30.rdResp_edirRam__00__1, m31.rdResp_edirRam__00__0,
    m8.rdResp_infoRam__00__15, m9.rdResp_infoRam__00__14,
    m10.rdResp_infoRam__00__13, m11.rdResp_infoRam__00__12,
    m12.rdResp_infoRam__00__11, m13.rdResp_infoRam__00__10,
    m14.rdResp_infoRam__00__9, m15.rdResp_infoRam__00__8,
    m16.rdResp_infoRam__00__7, m17.rdResp_infoRam__00__6,
    m18.rdResp_infoRam__00__5, m19.rdResp_infoRam__00__4,
    m20.rdResp_infoRam__00__3, m21.rdResp_infoRam__00__2,
    m22.rdResp_infoRam__00__1, m23.rdResp_infoRam__00__0, m7.enq_cp_2__00,
    m6.deq_cp_1__00, m157.repGetRq__00, m24.rdReq_edirRam__00__7,
    m25.rdReq_edirRam__00__6, m26.rdReq_edirRam__00__5,
    m27.rdReq_edirRam__00__4, m28.rdReq_edirRam__00__3,
    m29.rdReq_edirRam__00__2, m30.rdReq_edirRam__00__1,
    m31.rdReq_edirRam__00__0, m8.rdReq_infoRam__00__15,
    m9.rdReq_infoRam__00__14, m10.rdReq_infoRam__00__13,
    m11.rdReq_infoRam__00__12, m12.rdReq_infoRam__00__11,
    m13.rdReq_infoRam__00__10, m14.rdReq_infoRam__00__9,
    m15.rdReq_infoRam__00__8, m16.rdReq_infoRam__00__7,
    m17.rdReq_infoRam__00__6, m18.rdReq_infoRam__00__5,
    m19.rdReq_infoRam__00__4, m20.rdReq_infoRam__00__3,
    m21.rdReq_infoRam__00__2, m22.rdReq_infoRam__00__1,
    m23.rdReq_infoRam__00__0, m6.enq_cp_1__00);
    Module181 m181 <- mkModule181 (m53.wrReq_edirRam__000__3,
    m54.wrReq_edirRam__000__2, m55.wrReq_edirRam__000__1,
    m56.wrReq_edirRam__000__0, m57.wrReq_dataRam__000, m162.repAccess__000,
    m45.wrReq_infoRam__000__7, m46.wrReq_infoRam__000__6,
    m47.wrReq_infoRam__000__5, m48.wrReq_infoRam__000__4,
    m49.wrReq_infoRam__000__3, m50.wrReq_infoRam__000__2,
    m51.wrReq_infoRam__000__1, m52.wrReq_infoRam__000__0,
    m57.rdResp_dataRam__000, m44.deq_cp_2__000, m57.rdReq_dataRam__000,
    m162.repGetRs__000, m53.rdResp_edirRam__000__3,
    m54.rdResp_edirRam__000__2, m55.rdResp_edirRam__000__1,
    m56.rdResp_edirRam__000__0, m45.rdResp_infoRam__000__7,
    m46.rdResp_infoRam__000__6, m47.rdResp_infoRam__000__5,
    m48.rdResp_infoRam__000__4, m49.rdResp_infoRam__000__3,
    m50.rdResp_infoRam__000__2, m51.rdResp_infoRam__000__1,
    m52.rdResp_infoRam__000__0, m44.enq_cp_2__000, m43.deq_cp_1__000,
    m162.repGetRq__000, m53.rdReq_edirRam__000__3, m54.rdReq_edirRam__000__2,
    m55.rdReq_edirRam__000__1, m56.rdReq_edirRam__000__0,
    m45.rdReq_infoRam__000__7, m46.rdReq_infoRam__000__6,
    m47.rdReq_infoRam__000__5, m48.rdReq_infoRam__000__4,
    m49.rdReq_infoRam__000__3, m50.rdReq_infoRam__000__2,
    m51.rdReq_infoRam__000__1, m52.rdReq_infoRam__000__0, m43.enq_cp_1__000);

    Module182 m182 <- mkModule182 (m165.repAccess__0000,
    m74.wrReq_dataRam__0000, m70.wrReq_infoRam__0000__3,
    m71.wrReq_infoRam__0000__2, m72.wrReq_infoRam__0000__1,
    m73.wrReq_infoRam__0000__0, m74.rdResp_dataRam__0000, m69.deq_cp_2__0000,
    m74.rdReq_dataRam__0000, m165.repGetRs__0000,
    m70.rdResp_infoRam__0000__3, m71.rdResp_infoRam__0000__2,
    m72.rdResp_infoRam__0000__1, m73.rdResp_infoRam__0000__0,
    m69.enq_cp_2__0000, m68.deq_cp_1__0000, m165.repGetRq__0000,
    m70.rdReq_infoRam__0000__3, m71.rdReq_infoRam__0000__2,
    m72.rdReq_infoRam__0000__1, m73.rdReq_infoRam__0000__0,
    m68.enq_cp_1__0000);
    Module183 m183 <- mkModule183 (m168.repAccess__0001,
    m91.wrReq_dataRam__0001, m87.wrReq_infoRam__0001__3,
    m88.wrReq_infoRam__0001__2, m89.wrReq_infoRam__0001__1,
    m90.wrReq_infoRam__0001__0, m91.rdResp_dataRam__0001, m86.deq_cp_2__0001,
    m91.rdReq_dataRam__0001, m168.repGetRs__0001,
    m87.rdResp_infoRam__0001__3, m88.rdResp_infoRam__0001__2,
    m89.rdResp_infoRam__0001__1, m90.rdResp_infoRam__0001__0,
    m86.enq_cp_2__0001, m85.deq_cp_1__0001, m168.repGetRq__0001,
    m87.rdReq_infoRam__0001__3, m88.rdReq_infoRam__0001__2,
    m89.rdReq_infoRam__0001__1, m90.rdReq_infoRam__0001__0,
    m85.enq_cp_1__0001);
    Module184 m184 <- mkModule184 (m112.wrReq_edirRam__001__3,
    m113.wrReq_edirRam__001__2, m114.wrReq_edirRam__001__1,
    m115.wrReq_edirRam__001__0, m116.wrReq_dataRam__001, m173.repAccess__001,
    m104.wrReq_infoRam__001__7, m105.wrReq_infoRam__001__6,
    m106.wrReq_infoRam__001__5, m107.wrReq_infoRam__001__4,
    m108.wrReq_infoRam__001__3, m109.wrReq_infoRam__001__2,
    m110.wrReq_infoRam__001__1, m111.wrReq_infoRam__001__0,
    m116.rdResp_dataRam__001, m103.deq_cp_2__001, m116.rdReq_dataRam__001,
    m173.repGetRs__001, m112.rdResp_edirRam__001__3,
    m113.rdResp_edirRam__001__2, m114.rdResp_edirRam__001__1,
    m115.rdResp_edirRam__001__0, m104.rdResp_infoRam__001__7,
    m105.rdResp_infoRam__001__6, m106.rdResp_infoRam__001__5,
    m107.rdResp_infoRam__001__4, m108.rdResp_infoRam__001__3,
    m109.rdResp_infoRam__001__2, m110.rdResp_infoRam__001__1,
    m111.rdResp_infoRam__001__0, m103.enq_cp_2__001, m102.deq_cp_1__001,
    m173.repGetRq__001, m112.rdReq_edirRam__001__3,
    m113.rdReq_edirRam__001__2, m114.rdReq_edirRam__001__1,
    m115.rdReq_edirRam__001__0, m104.rdReq_infoRam__001__7,
    m105.rdReq_infoRam__001__6, m106.rdReq_infoRam__001__5,
    m107.rdReq_infoRam__001__4, m108.rdReq_infoRam__001__3,
    m109.rdReq_infoRam__001__2, m110.rdReq_infoRam__001__1,
    m111.rdReq_infoRam__001__0, m102.enq_cp_1__001);
    Module185 m185 <- mkModule185 (m176.repAccess__0010,
    m133.wrReq_dataRam__0010, m129.wrReq_infoRam__0010__3,
    m130.wrReq_infoRam__0010__2, m131.wrReq_infoRam__0010__1,
    m132.wrReq_infoRam__0010__0, m133.rdResp_dataRam__0010,
    m128.deq_cp_2__0010, m133.rdReq_dataRam__0010, m176.repGetRs__0010,
    m129.rdResp_infoRam__0010__3, m130.rdResp_infoRam__0010__2,
    m131.rdResp_infoRam__0010__1, m132.rdResp_infoRam__0010__0,
    m128.enq_cp_2__0010, m127.deq_cp_1__0010, m176.repGetRq__0010,
    m129.rdReq_infoRam__0010__3, m130.rdReq_infoRam__0010__2,
    m131.rdReq_infoRam__0010__1, m132.rdReq_infoRam__0010__0,
    m127.enq_cp_1__0010);
    Module186 m186 <- mkModule186 (m179.repAccess__0011,
    m150.wrReq_dataRam__0011, m146.wrReq_infoRam__0011__3,
    m147.wrReq_infoRam__0011__2, m148.wrReq_infoRam__0011__1,
    m149.wrReq_infoRam__0011__0, m150.rdResp_dataRam__0011,
    m145.deq_cp_2__0011, m150.rdReq_dataRam__0011, m179.repGetRs__0011,
    m146.rdResp_infoRam__0011__3, m147.rdResp_infoRam__0011__2,
    m148.rdResp_infoRam__0011__1, m149.rdResp_infoRam__0011__0,
    m145.enq_cp_2__0011, m144.deq_cp_1__0011, m179.repGetRq__0011,
    m146.rdReq_infoRam__0011__3, m147.rdReq_infoRam__0011__2,
    m148.rdReq_infoRam__0011__1, m149.rdReq_infoRam__0011__0,
    m144.enq_cp_1__0011);
    Module187 m187 <- mkModule187 (m180.cache__00__setVictimRq,
    m34.getULImm_00, m180.cache__00__getVictim, m34.transferUpDown_00,
    m156.broadcast_parentChildren00, m34.registerDL_00, m34.registerUL_00,
    m180.cache__00__getVictimCount, m34.getULCount_00,
    m156.makeEnq_parentChildren00, m180.cache__00__valueRsLineRq,
    m34.getMSHR_00, m5.deq_fifoL2E00, m5.enq_fifoL2E00,
    m180.cache__00__infoRsValueRq, m4.deq_fifoI2L00, m34.getRsReady_00,
    m34.releaseMSHR_00, m180.cache__00__releaseVictim, m34.getWait_00,
    m34.addRs_00, m34.getCRqSlot_00, m34.findUL_00, m4.enq_fifoI2L00,
    m180.cache__00__infoRq, m34.getPRqSlot_00, m3.deq_fifoInput00);
    Module188 m188 <- mkModule188 (m181.cache__000__setVictimRq,
    m59.getULImm_000, m181.cache__000__getVictim, m59.transferUpDown_000,
    m161.broadcast_parentChildren000, m59.registerDL_000, m59.registerUL_000,
    m181.cache__000__getVictimCount, m59.getULCount_000,
    m161.makeEnq_parentChildren000, m181.cache__000__valueRsLineRq,
    m59.getMSHR_000, m39.deq_fifoL2E000, m39.enq_fifoL2E000,
    m181.cache__000__infoRsValueRq, m38.deq_fifoI2L000, m59.getRsReady_000,
    m59.releaseMSHR_000, m181.cache__000__releaseVictim, m59.getWait_000,
    m59.addRs_000, m59.getCRqSlot_000, m59.findUL_000, m38.enq_fifoI2L000,
    m181.cache__000__infoRq, m59.getPRqSlot_000, m37.deq_fifoInput000);

    Module189 m189 <- mkModule189 (m182.cache__0000__setVictimRq,
    m76.getULImm_0000, m182.cache__0000__getVictim, m76.registerUL_0000,
    m182.cache__0000__getVictimCount, m76.getULCount_0000,
    m164.makeEnq_parentChildren0000, m182.cache__0000__valueRsLineRq,
    m76.getMSHR_0000, m62.deq_fifoL2E0000, m62.enq_fifoL2E0000,
    m182.cache__0000__infoRsValueRq, m61.deq_fifoI2L0000,
    m76.getRsReady_0000, m76.releaseMSHR_0000,
    m182.cache__0000__releaseVictim, m76.getWait_0000, m76.addRs_0000,
    m76.getCRqSlot_0000, m76.findUL_0000, m61.enq_fifoI2L0000,
    m182.cache__0000__infoRq, m76.getPRqSlot_0000, m60.deq_fifoInput0000);

    Module190 m190 <- mkModule190 (m183.cache__0001__setVictimRq,
    m93.getULImm_0001, m183.cache__0001__getVictim, m93.registerUL_0001,
    m183.cache__0001__getVictimCount, m93.getULCount_0001,
    m167.makeEnq_parentChildren0001, m183.cache__0001__valueRsLineRq,
    m93.getMSHR_0001, m79.deq_fifoL2E0001, m79.enq_fifoL2E0001,
    m183.cache__0001__infoRsValueRq, m78.deq_fifoI2L0001,
    m93.getRsReady_0001, m93.releaseMSHR_0001,
    m183.cache__0001__releaseVictim, m93.getWait_0001, m93.addRs_0001,
    m93.getCRqSlot_0001, m93.findUL_0001, m78.enq_fifoI2L0001,
    m183.cache__0001__infoRq, m93.getPRqSlot_0001, m77.deq_fifoInput0001);

    Module191 m191 <- mkModule191 (m184.cache__001__setVictimRq,
    m118.getULImm_001, m184.cache__001__getVictim, m118.transferUpDown_001,
    m172.broadcast_parentChildren001, m118.registerDL_001,
    m118.registerUL_001, m184.cache__001__getVictimCount,
    m118.getULCount_001, m172.makeEnq_parentChildren001,
    m184.cache__001__valueRsLineRq, m118.getMSHR_001, m98.deq_fifoL2E001,
    m98.enq_fifoL2E001, m184.cache__001__infoRsValueRq, m97.deq_fifoI2L001,
    m118.getRsReady_001, m118.releaseMSHR_001,
    m184.cache__001__releaseVictim, m118.getWait_001, m118.addRs_001,
    m118.getCRqSlot_001, m118.findUL_001, m97.enq_fifoI2L001,
    m184.cache__001__infoRq, m118.getPRqSlot_001, m96.deq_fifoInput001);

    Module192 m192 <- mkModule192 (m185.cache__0010__setVictimRq,
    m135.getULImm_0010, m185.cache__0010__getVictim, m135.registerUL_0010,
    m185.cache__0010__getVictimCount, m135.getULCount_0010,
    m175.makeEnq_parentChildren0010, m185.cache__0010__valueRsLineRq,
    m135.getMSHR_0010, m121.deq_fifoL2E0010, m121.enq_fifoL2E0010,
    m185.cache__0010__infoRsValueRq, m120.deq_fifoI2L0010,
    m135.getRsReady_0010, m135.releaseMSHR_0010,
    m185.cache__0010__releaseVictim, m135.getWait_0010, m135.addRs_0010,
    m135.getCRqSlot_0010, m135.findUL_0010, m120.enq_fifoI2L0010,
    m185.cache__0010__infoRq, m135.getPRqSlot_0010, m119.deq_fifoInput0010);

    Module193 m193 <- mkModule193 (m186.cache__0011__setVictimRq,
    m152.getULImm_0011, m186.cache__0011__getVictim, m152.registerUL_0011,
    m186.cache__0011__getVictimCount, m152.getULCount_0011,
    m178.makeEnq_parentChildren0011, m186.cache__0011__valueRsLineRq,
    m152.getMSHR_0011, m138.deq_fifoL2E0011, m138.enq_fifoL2E0011,
    m186.cache__0011__infoRsValueRq, m137.deq_fifoI2L0011,
    m152.getRsReady_0011, m152.releaseMSHR_0011,
    m186.cache__0011__releaseVictim, m152.getWait_0011, m152.addRs_0011,
    m152.getCRqSlot_0011, m152.findUL_0011, m137.enq_fifoI2L0011,
    m186.cache__0011__infoRq, m152.getPRqSlot_0011, m136.deq_fifoInput0011);

        //// Interface

    function MemRqRs getMemRqRs (function Action enq_rq (Struct1 _),
                                 function ActionValue#(Struct1) deq_rs ());
        return interface MemRqRs;
                   method mem_enq_rq = enq_rq;
                   method mem_deq_rs = deq_rs;
               endinterface;
    endfunction

    Vector#(L1Num, MemRqRs) _l1Ifc = newVector();
    _l1Ifc[0] = getMemRqRs(m66.enq_fifo000000, m67.deq_fifo000002);
    _l1Ifc[1] = getMemRqRs(m83.enq_fifo000100, m84.deq_fifo000102);
    _l1Ifc[2] = getMemRqRs(m125.enq_fifo001000, m126.deq_fifo001002);
    _l1Ifc[3] = getMemRqRs(m142.enq_fifo001100, m143.deq_fifo001102);
    interface l1Ifc = _l1Ifc;

    interface DMA llDma;
        method dma_rdReq = m32.rdReq_dataRam__00;
        method dma_wrReq = m32.wrReq_dataRam__00;
        method dma_rdResp = m32.rdResp_dataRam__00;
    endinterface

endmodule
