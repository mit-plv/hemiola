CCWrapper_L1LL.bsv