CC_L1LL2.bsv