import Vector::*;
import BuildVector::*;
import FIFO::*;
import FIFOF::*;
import RWBramCore::*;
import SpecialFIFOs::*;

typedef struct { Bool rl_valid; Bit#(2) rl_cmidx; Struct2 rl_msg; Bool rl_line_valid; Struct3 rl_line;  } Struct1 deriving(Eq, Bits);
typedef struct { Bit#(2) enq_type; Bit#(2) enq_ch_idx; Struct2 enq_msg;  } Struct10 deriving(Eq, Bits);
typedef struct { Bool r_ul_rsb; Struct2 r_ul_msg; Bit#(2) r_ul_rsbTo;  } Struct11 deriving(Eq, Bits);
typedef struct { Bool r_dl_rsb; Struct2 r_dl_msg; Bit#(4) r_dl_rss_from; Bit#(4) r_dl_rsbTo;  } Struct12 deriving(Eq, Bits);
typedef struct { Bit#(4) cs_inds; Struct2 cs_msg;  } Struct13 deriving(Eq, Bits);
typedef struct { Bit#(64) r_dl_addr; Bit#(2) r_dl_midx; Struct2 r_dl_msg;  } Struct14 deriving(Eq, Bits);
typedef struct { Bool valid; Struct9 data;  } Struct15 deriving(Eq, Bits);
typedef struct { Bit#(4) cidx; Struct2 msg;  } Struct16 deriving(Eq, Bits);
typedef struct { Bit#(64) r_dl_addr; Bit#(4) r_dl_rss_from;  } Struct17 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(3) victim_idx; Struct3 victim_line;  } Struct18 deriving(Eq, Bits);
typedef struct { Bit#(51) tag; Struct4 value;  } Struct19 deriving(Eq, Bits);
typedef struct { Bit#(6) id; Bool type_; Bit#(64) addr; Bit#(64) value;  } Struct2 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(4) tm_way; Struct4 tm_value;  } Struct20 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(14) addr; Bit#(64) datain;  } Struct21 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(10) addr; Struct19 datain;  } Struct22 deriving(Eq, Bits);
typedef struct { Bool rl_valid; Bit#(2) rl_cmidx; Struct2 rl_msg; Bool rl_line_valid; Struct24 rl_line;  } Struct23 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_hit; Bit#(3) info_way; Bool info_write; Struct4 info; Bool value_write; Bit#(64) value;  } Struct24 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(3) victim_idx; Struct24 victim_line;  } Struct25 deriving(Eq, Bits);
typedef struct { Bit#(53) tag; Struct4 value;  } Struct26 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(3) tm_way; Struct4 tm_value;  } Struct27 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(11) addr; Bit#(64) datain;  } Struct28 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(8) addr; Struct26 datain;  } Struct29 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_hit; Bit#(4) info_way; Bool info_write; Struct4 info; Bool value_write; Bit#(64) value;  } Struct3 deriving(Eq, Bits);
typedef struct { Bool rl_valid; Bit#(2) rl_cmidx; Struct2 rl_msg; Bool rl_line_valid; Struct31 rl_line;  } Struct30 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_hit; Bit#(2) info_way; Bool info_write; Struct4 info; Bool value_write; Bit#(64) value;  } Struct31 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(2) victim_idx; Struct31 victim_line;  } Struct32 deriving(Eq, Bits);
typedef struct { Bit#(55) tag; Struct4 value;  } Struct33 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(2) tm_way; Struct4 tm_value;  } Struct34 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(8) addr; Bit#(64) datain;  } Struct35 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(6) addr; Struct33 datain;  } Struct36 deriving(Eq, Bits);
typedef struct { Bool mesi_owned; Bit#(3) mesi_status; Bit#(3) mesi_dir_st; Bit#(4) mesi_dir_sharers;  } Struct4 deriving(Eq, Bits);
typedef struct { Bool wl_valid; Bool wl_write_rq;  } Struct5 deriving(Eq, Bits);
typedef struct { Bool valid; Struct7 data;  } Struct6 deriving(Eq, Bits);
typedef struct { Bool dl_valid; Bool dl_rsb; Struct2 dl_msg; Bit#(4) dl_rss_from; Bit#(4) dl_rss_recv; Vector#(4, Struct2) dl_rss; Bit#(4) dl_rsbTo;  } Struct7 deriving(Eq, Bits);
typedef struct { Bit#(3) dir_st; Bit#(2) dir_excl; Bit#(4) dir_sharers;  } Struct8 deriving(Eq, Bits);
typedef struct { Bool ul_valid; Bool ul_rsb; Struct2 ul_msg; Bit#(2) ul_rsbTo;  } Struct9 deriving(Eq, Bits);

interface Module1;
    method Action putRq_infoRam_00_15 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_15 ();

endinterface

module mkModule1 (Module1);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_15 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_15 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module2;
    method Action putRq_infoRam_00_14 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_14 ();

endinterface

module mkModule2 (Module2);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_14 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_14 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module3;
    method Action putRq_infoRam_00_13 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_13 ();

endinterface

module mkModule3 (Module3);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_13 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_13 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module4;
    method Action putRq_infoRam_00_12 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_12 ();

endinterface

module mkModule4 (Module4);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_12 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_12 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module5;
    method Action putRq_infoRam_00_11 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_11 ();

endinterface

module mkModule5 (Module5);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_11 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_11 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module6;
    method Action putRq_infoRam_00_10 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_10 ();

endinterface

module mkModule6 (Module6);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_10 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_10 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module7;
    method Action putRq_infoRam_00_9 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_9 ();

endinterface

module mkModule7 (Module7);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_9 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_9 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module8;
    method Action putRq_infoRam_00_8 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_8 ();

endinterface

module mkModule8 (Module8);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_8 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_8 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module9;
    method Action putRq_infoRam_00_7 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_7 ();

endinterface

module mkModule9 (Module9);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_7 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_7 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module10;
    method Action putRq_infoRam_00_6 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_6 ();

endinterface

module mkModule10 (Module10);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_6 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_6 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module11;
    method Action putRq_infoRam_00_5 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_5 ();

endinterface

module mkModule11 (Module11);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_5 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_5 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module12;
    method Action putRq_infoRam_00_4 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_4 ();

endinterface

module mkModule12 (Module12);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_4 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_4 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module13;
    method Action putRq_infoRam_00_3 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_3 ();

endinterface

module mkModule13 (Module13);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_3 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module14;
    method Action putRq_infoRam_00_2 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_2 ();

endinterface

module mkModule14 (Module14);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_2 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module15;
    method Action putRq_infoRam_00_1 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_1 ();

endinterface

module mkModule15 (Module15);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_1 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module16;
    method Action putRq_infoRam_00_0 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_0 ();

endinterface

module mkModule16 (Module16);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_0 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module17;
    method Action putRq_dataRam_00 (Struct21 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_00 ();

endinterface

module mkModule17 (Module17);
    RWBramCore#(Bit#(14), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_00 (Struct21 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_00 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module18;
    method ActionValue#(Bool) upLockable00 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable00 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet00 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet00 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull00 ();
    method Action registerUL00 (Struct11 x_0);
    method Action releaseUL00 (Bit#(64) x_0);
    method Action registerDL00 (Struct12 x_0);
    method Action releaseDL00 (Bit#(64) x_0);
    method Action transferUpDown00 (Struct17 x_0);
    method Action addRs00 (Struct14 x_0);

endinterface

module mkModule18 (Module18);
    Reg#(Vector#(8, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(8, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable00 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(3))'(3'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h3)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h4)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h5)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h6)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h7)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))))))))))));
        Bool x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable00 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(3))'(3'h1)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h2)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h3)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h4)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h5)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h6)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h7)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))))))))))));
        Bool x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h4)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h5)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h6)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h7)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet00 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h0)]}) :
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h1)]}) :
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h2)]}) :
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h3)]}) :
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h4)]}) :
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h5)]}) :
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h6)]}) :
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h7)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet00 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h0)]}) :
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h1)]}) :
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h2)]}) :
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h3)]}) :
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h4)]}) :
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h5)]}) :
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h6)]}) :
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h7)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull00 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h0)]}) :
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h1)]}) :
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h2)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h2)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h2)]}) :
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h3)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h3)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h3)]}) :
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h4)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h4)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h4)]}) :
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h5)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h5)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h5)]}) :
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h6)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h6)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h6)]}) :
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_valid) &&
        ((((x_1)[(Bit#(3))'(3'h7)]).dl_rss_recv) ==
        (((x_1)[(Bit#(3))'(3'h7)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h7)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))))))))))));

        return x_2;
    endmethod

    method Action registerUL00 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(3) x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).ul_valid) ?
        ((Bit#(3))'(3'h0)) : ((! (((x_1)[(Bit#(3))'(3'h1)]).ul_valid) ?
        ((Bit#(3))'(3'h1)) : ((! (((x_1)[(Bit#(3))'(3'h2)]).ul_valid) ?
        ((Bit#(3))'(3'h2)) : ((! (((x_1)[(Bit#(3))'(3'h3)]).ul_valid) ?
        ((Bit#(3))'(3'h3)) : ((! (((x_1)[(Bit#(3))'(3'h4)]).ul_valid) ?
        ((Bit#(3))'(3'h4)) : ((! (((x_1)[(Bit#(3))'(3'h5)]).ul_valid) ?
        ((Bit#(3))'(3'h5)) : ((! (((x_1)[(Bit#(3))'(3'h6)]).ul_valid) ?
        ((Bit#(3))'(3'h6)) : ((! (((x_1)[(Bit#(3))'(3'h7)]).ul_valid) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL00 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL00 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(3) x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).dl_valid) ?
        ((Bit#(3))'(3'h0)) : ((! (((x_1)[(Bit#(3))'(3'h1)]).dl_valid) ?
        ((Bit#(3))'(3'h1)) : ((! (((x_1)[(Bit#(3))'(3'h2)]).dl_valid) ?
        ((Bit#(3))'(3'h2)) : ((! (((x_1)[(Bit#(3))'(3'h3)]).dl_valid) ?
        ((Bit#(3))'(3'h3)) : ((! (((x_1)[(Bit#(3))'(3'h4)]).dl_valid) ?
        ((Bit#(3))'(3'h4)) : ((! (((x_1)[(Bit#(3))'(3'h5)]).dl_valid) ?
        ((Bit#(3))'(3'h5)) : ((! (((x_1)[(Bit#(3))'(3'h6)]).dl_valid) ?
        ((Bit#(3))'(3'h6)) : ((! (((x_1)[(Bit#(3))'(3'h7)]).dl_valid) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL00 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown00 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(3) x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(3) x_6 = ((! (((x_5)[(Bit#(3))'(3'h0)]).dl_valid) ?
        ((Bit#(3))'(3'h0)) : ((! (((x_5)[(Bit#(3))'(3'h1)]).dl_valid) ?
        ((Bit#(3))'(3'h1)) : ((! (((x_5)[(Bit#(3))'(3'h2)]).dl_valid) ?
        ((Bit#(3))'(3'h2)) : ((! (((x_5)[(Bit#(3))'(3'h3)]).dl_valid) ?
        ((Bit#(3))'(3'h3)) : ((! (((x_5)[(Bit#(3))'(3'h4)]).dl_valid) ?
        ((Bit#(3))'(3'h4)) : ((! (((x_5)[(Bit#(3))'(3'h5)]).dl_valid) ?
        ((Bit#(3))'(3'h5)) : ((! (((x_5)[(Bit#(3))'(3'h6)]).dl_valid) ?
        ((Bit#(3))'(3'h6)) : ((! (((x_5)[(Bit#(3))'(3'h7)]).dl_valid) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs00 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        Struct6 x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h0)]}) :
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h1)]}) :
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h2)]}) :
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h3)]}) :
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h4)]}) :
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h5)]}) :
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h6)]}) :
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h7)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))))))))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module19;
    method Action putRq_infoRam_000_7 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_7 ();

endinterface

module mkModule19 (Module19);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_7 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_7 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module20;
    method Action putRq_infoRam_000_6 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_6 ();

endinterface

module mkModule20 (Module20);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_6 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_6 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module21;
    method Action putRq_infoRam_000_5 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_5 ();

endinterface

module mkModule21 (Module21);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_5 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_5 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module22;
    method Action putRq_infoRam_000_4 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_4 ();

endinterface

module mkModule22 (Module22);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_4 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_4 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module23;
    method Action putRq_infoRam_000_3 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_3 ();

endinterface

module mkModule23 (Module23);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_3 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module24;
    method Action putRq_infoRam_000_2 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_2 ();

endinterface

module mkModule24 (Module24);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_2 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module25;
    method Action putRq_infoRam_000_1 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_1 ();

endinterface

module mkModule25 (Module25);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_1 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module26;
    method Action putRq_infoRam_000_0 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_0 ();

endinterface

module mkModule26 (Module26);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_0 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module27;
    method Action putRq_dataRam_000 (Struct28 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_000 ();

endinterface

module mkModule27 (Module27);
    RWBramCore#(Bit#(11), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_000 (Struct28 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_000 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module28;
    method ActionValue#(Bool) upLockable000 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable000 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet000 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet000 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull000 ();
    method Action registerUL000 (Struct11 x_0);
    method Action releaseUL000 (Bit#(64) x_0);
    method Action registerDL000 (Struct12 x_0);
    method Action releaseDL000 (Bit#(64) x_0);
    method Action transferUpDown000 (Struct17 x_0);
    method Action addRs000 (Struct14 x_0);

endinterface

module mkModule28 (Module28);
    Reg#(Vector#(8, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable000 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(3))'(3'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h3)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h4)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h5)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h6)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h7)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))))))))))));
        Bool x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable000 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet000 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h0)]}) :
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h1)]}) :
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h2)]}) :
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h3)]}) :
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h4)]}) :
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h5)]}) :
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h6)]}) :
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h7)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet000 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull000 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h2)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h2)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h3)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h3)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))));

        return x_2;
    endmethod

    method Action registerUL000 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(3) x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).ul_valid) ?
        ((Bit#(3))'(3'h0)) : ((! (((x_1)[(Bit#(3))'(3'h1)]).ul_valid) ?
        ((Bit#(3))'(3'h1)) : ((! (((x_1)[(Bit#(3))'(3'h2)]).ul_valid) ?
        ((Bit#(3))'(3'h2)) : ((! (((x_1)[(Bit#(3))'(3'h3)]).ul_valid) ?
        ((Bit#(3))'(3'h3)) : ((! (((x_1)[(Bit#(3))'(3'h4)]).ul_valid) ?
        ((Bit#(3))'(3'h4)) : ((! (((x_1)[(Bit#(3))'(3'h5)]).ul_valid) ?
        ((Bit#(3))'(3'h5)) : ((! (((x_1)[(Bit#(3))'(3'h6)]).ul_valid) ?
        ((Bit#(3))'(3'h6)) : ((! (((x_1)[(Bit#(3))'(3'h7)]).ul_valid) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL000 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL000 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).dl_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).dl_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).dl_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).dl_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL000 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown000 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(3) x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(2) x_6 = ((! (((x_5)[(Bit#(2))'(2'h0)]).dl_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_5)[(Bit#(2))'(2'h1)]).dl_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_5)[(Bit#(2))'(2'h2)]).dl_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_5)[(Bit#(2))'(2'h3)]).dl_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs000 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct6 x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module29;
    method Action enq_fifo0000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0000 ();

endinterface

module mkModule29 (Module29);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo0000 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0000 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module30;
    method Action enq_fifo0001 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0001 ();

endinterface

module mkModule30 (Module30);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo0001 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0001 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module31;
    method Action enq_fifo0002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0002 ();

endinterface

module mkModule31 (Module31);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo0002 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0002 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module32;
    method Action putRq_infoRam_0000_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0000_3 ();

endinterface

module mkModule32 (Module32);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0000_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0000_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module33;
    method Action putRq_infoRam_0000_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0000_2 ();

endinterface

module mkModule33 (Module33);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0000_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0000_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module34;
    method Action putRq_infoRam_0000_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0000_1 ();

endinterface

module mkModule34 (Module34);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0000_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0000_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module35;
    method Action putRq_infoRam_0000_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0000_0 ();

endinterface

module mkModule35 (Module35);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0000_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0000_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module36;
    method Action putRq_dataRam_0000 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0000 ();

endinterface

module mkModule36 (Module36);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0000 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0000 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module37;
    method ActionValue#(Bool) upLockable0000 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0000 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0000 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0000 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0000 ();
    method Action registerUL0000 (Struct11 x_0);
    method Action releaseUL0000 (Bit#(64) x_0);
    method Action registerDL0000 (Struct12 x_0);
    method Action releaseDL0000 (Bit#(64) x_0);
    method Action transferUpDown0000 (Struct17 x_0);
    method Action addRs0000 (Struct14 x_0);

endinterface

module mkModule37 (Module37);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0000 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0000 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0000 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0000 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0000 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0000 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0000 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0000 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0000 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0000 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0000 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module38;
    method Action enq_fifo00000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00000 ();

endinterface

module mkModule38 (Module38);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00000 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00000 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module39;
    method Action enq_fifo00001 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00001 ();

endinterface

module mkModule39 (Module39);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00001 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00001 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module40;
    method Action enq_fifo00002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00002 ();

endinterface

module mkModule40 (Module40);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00002 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00002 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module41;
    method Action enq_fifo000000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000000 ();

endinterface

module mkModule41 (Module41);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000000 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000000 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module42;
    method Action enq_fifo000002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000002 ();

endinterface

module mkModule42 (Module42);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000002 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000002 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module43;
    method Action putRq_infoRam_0001_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0001_3 ();

endinterface

module mkModule43 (Module43);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0001_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0001_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module44;
    method Action putRq_infoRam_0001_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0001_2 ();

endinterface

module mkModule44 (Module44);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0001_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0001_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module45;
    method Action putRq_infoRam_0001_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0001_1 ();

endinterface

module mkModule45 (Module45);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0001_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0001_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module46;
    method Action putRq_infoRam_0001_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0001_0 ();

endinterface

module mkModule46 (Module46);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0001_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0001_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module47;
    method Action putRq_dataRam_0001 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0001 ();

endinterface

module mkModule47 (Module47);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0001 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0001 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module48;
    method ActionValue#(Bool) upLockable0001 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0001 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0001 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0001 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0001 ();
    method Action registerUL0001 (Struct11 x_0);
    method Action releaseUL0001 (Bit#(64) x_0);
    method Action registerDL0001 (Struct12 x_0);
    method Action releaseDL0001 (Bit#(64) x_0);
    method Action transferUpDown0001 (Struct17 x_0);
    method Action addRs0001 (Struct14 x_0);

endinterface

module mkModule48 (Module48);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0001 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0001 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0001 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0001 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0001 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0001 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0001 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0001 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0001 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0001 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0001 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module49;
    method Action enq_fifo00010 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00010 ();

endinterface

module mkModule49 (Module49);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00010 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00010 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module50;
    method Action enq_fifo00011 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00011 ();

endinterface

module mkModule50 (Module50);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00011 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00011 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module51;
    method Action enq_fifo00012 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00012 ();

endinterface

module mkModule51 (Module51);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00012 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00012 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module52;
    method Action enq_fifo000100 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000100 ();

endinterface

module mkModule52 (Module52);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000100 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000100 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module53;
    method Action enq_fifo000102 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000102 ();

endinterface

module mkModule53 (Module53);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000102 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000102 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module54;
    method Action putRq_infoRam_0002_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0002_3 ();

endinterface

module mkModule54 (Module54);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0002_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0002_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module55;
    method Action putRq_infoRam_0002_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0002_2 ();

endinterface

module mkModule55 (Module55);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0002_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0002_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module56;
    method Action putRq_infoRam_0002_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0002_1 ();

endinterface

module mkModule56 (Module56);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0002_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0002_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module57;
    method Action putRq_infoRam_0002_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0002_0 ();

endinterface

module mkModule57 (Module57);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0002_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0002_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module58;
    method Action putRq_dataRam_0002 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0002 ();

endinterface

module mkModule58 (Module58);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0002 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0002 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module59;
    method ActionValue#(Bool) upLockable0002 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0002 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0002 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0002 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0002 ();
    method Action registerUL0002 (Struct11 x_0);
    method Action releaseUL0002 (Bit#(64) x_0);
    method Action registerDL0002 (Struct12 x_0);
    method Action releaseDL0002 (Bit#(64) x_0);
    method Action transferUpDown0002 (Struct17 x_0);
    method Action addRs0002 (Struct14 x_0);

endinterface

module mkModule59 (Module59);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0002 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0002 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0002 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0002 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0002 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0002 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0002 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0002 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0002 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0002 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0002 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module60;
    method Action enq_fifo00020 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00020 ();

endinterface

module mkModule60 (Module60);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00020 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00020 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module61;
    method Action enq_fifo00021 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00021 ();

endinterface

module mkModule61 (Module61);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00021 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00021 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module62;
    method Action enq_fifo00022 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00022 ();

endinterface

module mkModule62 (Module62);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00022 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00022 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module63;
    method Action enq_fifo000200 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000200 ();

endinterface

module mkModule63 (Module63);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000200 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000200 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module64;
    method Action enq_fifo000202 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000202 ();

endinterface

module mkModule64 (Module64);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000202 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000202 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module65;
    method Action putRq_infoRam_0003_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0003_3 ();

endinterface

module mkModule65 (Module65);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0003_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0003_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module66;
    method Action putRq_infoRam_0003_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0003_2 ();

endinterface

module mkModule66 (Module66);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0003_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0003_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module67;
    method Action putRq_infoRam_0003_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0003_1 ();

endinterface

module mkModule67 (Module67);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0003_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0003_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module68;
    method Action putRq_infoRam_0003_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0003_0 ();

endinterface

module mkModule68 (Module68);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0003_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0003_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module69;
    method Action putRq_dataRam_0003 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0003 ();

endinterface

module mkModule69 (Module69);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0003 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0003 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module70;
    method ActionValue#(Bool) upLockable0003 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0003 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0003 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0003 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0003 ();
    method Action registerUL0003 (Struct11 x_0);
    method Action releaseUL0003 (Bit#(64) x_0);
    method Action registerDL0003 (Struct12 x_0);
    method Action releaseDL0003 (Bit#(64) x_0);
    method Action transferUpDown0003 (Struct17 x_0);
    method Action addRs0003 (Struct14 x_0);

endinterface

module mkModule70 (Module70);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0003 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0003 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0003 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0003 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0003 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0003 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0003 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0003 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0003 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0003 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0003 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module71;
    method Action enq_fifo00030 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00030 ();

endinterface

module mkModule71 (Module71);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00030 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00030 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module72;
    method Action enq_fifo00031 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00031 ();

endinterface

module mkModule72 (Module72);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00031 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00031 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module73;
    method Action enq_fifo00032 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00032 ();

endinterface

module mkModule73 (Module73);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00032 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00032 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module74;
    method Action enq_fifo000300 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000300 ();

endinterface

module mkModule74 (Module74);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000300 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000300 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module75;
    method Action enq_fifo000302 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo000302 ();

endinterface

module mkModule75 (Module75);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo000302 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo000302 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module76;
    method Action putRq_infoRam_001_7 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_7 ();

endinterface

module mkModule76 (Module76);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_7 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_7 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module77;
    method Action putRq_infoRam_001_6 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_6 ();

endinterface

module mkModule77 (Module77);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_6 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_6 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module78;
    method Action putRq_infoRam_001_5 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_5 ();

endinterface

module mkModule78 (Module78);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_5 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_5 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module79;
    method Action putRq_infoRam_001_4 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_4 ();

endinterface

module mkModule79 (Module79);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_4 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_4 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module80;
    method Action putRq_infoRam_001_3 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_3 ();

endinterface

module mkModule80 (Module80);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_3 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module81;
    method Action putRq_infoRam_001_2 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_2 ();

endinterface

module mkModule81 (Module81);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_2 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module82;
    method Action putRq_infoRam_001_1 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_1 ();

endinterface

module mkModule82 (Module82);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_1 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module83;
    method Action putRq_infoRam_001_0 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_0 ();

endinterface

module mkModule83 (Module83);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_0 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module84;
    method Action putRq_dataRam_001 (Struct28 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_001 ();

endinterface

module mkModule84 (Module84);
    RWBramCore#(Bit#(11), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_001 (Struct28 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_001 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module85;
    method ActionValue#(Bool) upLockable001 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable001 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet001 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet001 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull001 ();
    method Action registerUL001 (Struct11 x_0);
    method Action releaseUL001 (Bit#(64) x_0);
    method Action registerDL001 (Struct12 x_0);
    method Action releaseDL001 (Bit#(64) x_0);
    method Action transferUpDown001 (Struct17 x_0);
    method Action addRs001 (Struct14 x_0);

endinterface

module mkModule85 (Module85);
    Reg#(Vector#(8, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable001 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(3))'(3'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h3)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h4)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h5)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h6)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(3))'(3'h7)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))))))))))));
        Bool x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable001 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet001 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h0)]}) :
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h1)]}) :
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h2)]}) :
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h3)]}) :
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h4)]}) :
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h5)]}) :
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h6)]}) :
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(3))'(3'h7)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet001 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull001 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h2)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h2)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h3)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h3)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))));

        return x_2;
    endmethod

    method Action registerUL001 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(3) x_2 = ((! (((x_1)[(Bit#(3))'(3'h0)]).ul_valid) ?
        ((Bit#(3))'(3'h0)) : ((! (((x_1)[(Bit#(3))'(3'h1)]).ul_valid) ?
        ((Bit#(3))'(3'h1)) : ((! (((x_1)[(Bit#(3))'(3'h2)]).ul_valid) ?
        ((Bit#(3))'(3'h2)) : ((! (((x_1)[(Bit#(3))'(3'h3)]).ul_valid) ?
        ((Bit#(3))'(3'h3)) : ((! (((x_1)[(Bit#(3))'(3'h4)]).ul_valid) ?
        ((Bit#(3))'(3'h4)) : ((! (((x_1)[(Bit#(3))'(3'h5)]).ul_valid) ?
        ((Bit#(3))'(3'h5)) : ((! (((x_1)[(Bit#(3))'(3'h6)]).ul_valid) ?
        ((Bit#(3))'(3'h6)) : ((! (((x_1)[(Bit#(3))'(3'h7)]).ul_valid) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL001 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(3) x_2 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL001 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).dl_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).dl_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).dl_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).dl_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL001 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown001 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(3) x_3 = (((((x_1)[(Bit#(3))'(3'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h0)) : (((((x_1)[(Bit#(3))'(3'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h1)) : (((((x_1)[(Bit#(3))'(3'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h2)) : (((((x_1)[(Bit#(3))'(3'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h3)) : (((((x_1)[(Bit#(3))'(3'h4)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h4)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h4)) : (((((x_1)[(Bit#(3))'(3'h5)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h5)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h5)) : (((((x_1)[(Bit#(3))'(3'h6)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h6)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h6)) : (((((x_1)[(Bit#(3))'(3'h7)]).ul_valid) &&
        (((((x_1)[(Bit#(3))'(3'h7)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h0))))))))))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(2) x_6 = ((! (((x_5)[(Bit#(2))'(2'h0)]).dl_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_5)[(Bit#(2))'(2'h1)]).dl_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_5)[(Bit#(2))'(2'h2)]).dl_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_5)[(Bit#(2))'(2'h3)]).dl_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs001 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct6 x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module86;
    method Action enq_fifo0010 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0010 ();

endinterface

module mkModule86 (Module86);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo0010 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0010 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module87;
    method Action enq_fifo0011 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0011 ();

endinterface

module mkModule87 (Module87);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo0011 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0011 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module88;
    method Action enq_fifo0012 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0012 ();

endinterface

module mkModule88 (Module88);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo0012 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0012 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module89;
    method Action putRq_infoRam_0010_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0010_3 ();

endinterface

module mkModule89 (Module89);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0010_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0010_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module90;
    method Action putRq_infoRam_0010_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0010_2 ();

endinterface

module mkModule90 (Module90);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0010_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0010_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module91;
    method Action putRq_infoRam_0010_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0010_1 ();

endinterface

module mkModule91 (Module91);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0010_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0010_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module92;
    method Action putRq_infoRam_0010_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0010_0 ();

endinterface

module mkModule92 (Module92);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0010_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0010_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module93;
    method Action putRq_dataRam_0010 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0010 ();

endinterface

module mkModule93 (Module93);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0010 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0010 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module94;
    method ActionValue#(Bool) upLockable0010 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0010 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0010 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0010 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0010 ();
    method Action registerUL0010 (Struct11 x_0);
    method Action releaseUL0010 (Bit#(64) x_0);
    method Action registerDL0010 (Struct12 x_0);
    method Action releaseDL0010 (Bit#(64) x_0);
    method Action transferUpDown0010 (Struct17 x_0);
    method Action addRs0010 (Struct14 x_0);

endinterface

module mkModule94 (Module94);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0010 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0010 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0010 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0010 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0010 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0010 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0010 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0010 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0010 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0010 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0010 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module95;
    method Action enq_fifo00100 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00100 ();

endinterface

module mkModule95 (Module95);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00100 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00100 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module96;
    method Action enq_fifo00101 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00101 ();

endinterface

module mkModule96 (Module96);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00101 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00101 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module97;
    method Action enq_fifo00102 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00102 ();

endinterface

module mkModule97 (Module97);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00102 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00102 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module98;
    method Action enq_fifo001000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001000 ();

endinterface

module mkModule98 (Module98);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001000 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001000 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module99;
    method Action enq_fifo001002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001002 ();

endinterface

module mkModule99 (Module99);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001002 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001002 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module100;
    method Action putRq_infoRam_0011_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0011_3 ();

endinterface

module mkModule100 (Module100);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0011_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0011_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module101;
    method Action putRq_infoRam_0011_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0011_2 ();

endinterface

module mkModule101 (Module101);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0011_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0011_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module102;
    method Action putRq_infoRam_0011_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0011_1 ();

endinterface

module mkModule102 (Module102);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0011_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0011_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module103;
    method Action putRq_infoRam_0011_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0011_0 ();

endinterface

module mkModule103 (Module103);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0011_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0011_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module104;
    method Action putRq_dataRam_0011 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0011 ();

endinterface

module mkModule104 (Module104);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0011 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0011 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module105;
    method ActionValue#(Bool) upLockable0011 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0011 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0011 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0011 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0011 ();
    method Action registerUL0011 (Struct11 x_0);
    method Action releaseUL0011 (Bit#(64) x_0);
    method Action registerDL0011 (Struct12 x_0);
    method Action releaseDL0011 (Bit#(64) x_0);
    method Action transferUpDown0011 (Struct17 x_0);
    method Action addRs0011 (Struct14 x_0);

endinterface

module mkModule105 (Module105);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0011 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0011 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0011 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0011 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0011 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0011 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0011 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0011 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0011 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0011 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0011 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module106;
    method Action enq_fifo00110 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00110 ();

endinterface

module mkModule106 (Module106);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00110 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00110 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module107;
    method Action enq_fifo00111 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00111 ();

endinterface

module mkModule107 (Module107);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00111 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00111 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module108;
    method Action enq_fifo00112 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00112 ();

endinterface

module mkModule108 (Module108);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00112 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00112 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module109;
    method Action enq_fifo001100 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001100 ();

endinterface

module mkModule109 (Module109);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001100 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001100 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module110;
    method Action enq_fifo001102 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001102 ();

endinterface

module mkModule110 (Module110);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001102 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001102 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module111;
    method Action putRq_infoRam_0012_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0012_3 ();

endinterface

module mkModule111 (Module111);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0012_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0012_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module112;
    method Action putRq_infoRam_0012_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0012_2 ();

endinterface

module mkModule112 (Module112);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0012_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0012_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module113;
    method Action putRq_infoRam_0012_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0012_1 ();

endinterface

module mkModule113 (Module113);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0012_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0012_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module114;
    method Action putRq_infoRam_0012_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0012_0 ();

endinterface

module mkModule114 (Module114);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0012_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0012_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module115;
    method Action putRq_dataRam_0012 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0012 ();

endinterface

module mkModule115 (Module115);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0012 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0012 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module116;
    method ActionValue#(Bool) upLockable0012 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0012 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0012 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0012 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0012 ();
    method Action registerUL0012 (Struct11 x_0);
    method Action releaseUL0012 (Bit#(64) x_0);
    method Action registerDL0012 (Struct12 x_0);
    method Action releaseDL0012 (Bit#(64) x_0);
    method Action transferUpDown0012 (Struct17 x_0);
    method Action addRs0012 (Struct14 x_0);

endinterface

module mkModule116 (Module116);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0012 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0012 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0012 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0012 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0012 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0012 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0012 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0012 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0012 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0012 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0012 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module117;
    method Action enq_fifo00120 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00120 ();

endinterface

module mkModule117 (Module117);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00120 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00120 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module118;
    method Action enq_fifo00121 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00121 ();

endinterface

module mkModule118 (Module118);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00121 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00121 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module119;
    method Action enq_fifo00122 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00122 ();

endinterface

module mkModule119 (Module119);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00122 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00122 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module120;
    method Action enq_fifo001200 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001200 ();

endinterface

module mkModule120 (Module120);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001200 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001200 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module121;
    method Action enq_fifo001202 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001202 ();

endinterface

module mkModule121 (Module121);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001202 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001202 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module122;
    method Action putRq_infoRam_0013_3 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0013_3 ();

endinterface

module mkModule122 (Module122);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0013_3 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0013_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module123;
    method Action putRq_infoRam_0013_2 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0013_2 ();

endinterface

module mkModule123 (Module123);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0013_2 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0013_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module124;
    method Action putRq_infoRam_0013_1 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0013_1 ();

endinterface

module mkModule124 (Module124);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0013_1 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0013_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module125;
    method Action putRq_infoRam_0013_0 (Struct36 x_0);
    method ActionValue#(Struct33) getRs_infoRam_0013_0 ();

endinterface

module mkModule125 (Module125);
    RWBramCore#(Bit#(6), Struct33) bram <- mkRWBramCore();

    method Action putRq_infoRam_0013_0 (Struct36 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct33) getRs_infoRam_0013_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module126;
    method Action putRq_dataRam_0013 (Struct35 x_0);
    method ActionValue#(Bit#(64)) getRs_dataRam_0013 ();

endinterface

module mkModule126 (Module126);
    RWBramCore#(Bit#(8), Bit#(64)) bram <- mkRWBramCore();

    method Action putRq_dataRam_0013 (Struct35 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Bit#(64)) getRs_dataRam_0013 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module127;
    method ActionValue#(Bool) upLockable0013 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable0013 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet0013 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet0013 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull0013 ();
    method Action registerUL0013 (Struct11 x_0);
    method Action releaseUL0013 (Bit#(64) x_0);
    method Action registerDL0013 (Struct12 x_0);
    method Action releaseDL0013 (Bit#(64) x_0);
    method Action transferUpDown0013 (Struct17 x_0);
    method Action addRs0013 (Struct14 x_0);

endinterface

module mkModule127 (Module127);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable0013 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable0013 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet0013 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet0013 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull0013 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL0013 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL0013 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL0013 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL0013 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown0013 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs0013 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module128;
    method Action enq_fifo00130 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00130 ();

endinterface

module mkModule128 (Module128);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00130 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00130 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module129;
    method Action enq_fifo00131 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00131 ();

endinterface

module mkModule129 (Module129);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00131 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00131 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module130;
    method Action enq_fifo00132 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00132 ();

endinterface

module mkModule130 (Module130);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo00132 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00132 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module131;
    method Action enq_fifo001300 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001300 ();

endinterface

module mkModule131 (Module131);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001300 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001300 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module132;
    method Action enq_fifo001302 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo001302 ();

endinterface

module mkModule132 (Module132);
    FIFOF#(Struct2) pff <- mkFIFOF();

    method Action enq_fifo001302 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo001302 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module133;
    method Action cache_00_readRq (Bit#(64) x_0);
    method ActionValue#(Struct3) cache_00_readRs ();
    method Action cache_00_writeRq (Struct3 x_0);
    method ActionValue#(Struct3) cache_00_writeRs ();
    method ActionValue#(Bool) cache_00_hasVictimSlot ();
    method ActionValue#(Struct3) cache_00_getVictim ();
    method Action cache_00_removeVictim (Bit#(64) x_0);

endinterface


module mkModule133#(function Action putRq_infoRam_00_15(Struct22 _),
  function Action putRq_infoRam_00_14(Struct22 _),
  function Action putRq_infoRam_00_13(Struct22 _),
  function Action putRq_infoRam_00_12(Struct22 _),
  function Action putRq_infoRam_00_11(Struct22 _),
  function Action putRq_infoRam_00_10(Struct22 _),
  function Action putRq_infoRam_00_9(Struct22 _),
  function Action putRq_infoRam_00_8(Struct22 _),
  function Action putRq_infoRam_00_7(Struct22 _),
  function Action putRq_infoRam_00_6(Struct22 _),
  function Action putRq_infoRam_00_5(Struct22 _),
  function Action putRq_infoRam_00_4(Struct22 _),
  function Action putRq_infoRam_00_3(Struct22 _),
  function Action putRq_infoRam_00_2(Struct22 _),
  function Action putRq_infoRam_00_1(Struct22 _),
  function Action putRq_infoRam_00_0(Struct22 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_00(),
  function Action putRq_dataRam_00(Struct21 _),
  function ActionValue#(Struct19) getRs_infoRam_00_15(),
  function ActionValue#(Struct19) getRs_infoRam_00_14(),
  function ActionValue#(Struct19) getRs_infoRam_00_13(),
  function ActionValue#(Struct19) getRs_infoRam_00_12(),
  function ActionValue#(Struct19) getRs_infoRam_00_11(),
  function ActionValue#(Struct19) getRs_infoRam_00_10(),
  function ActionValue#(Struct19) getRs_infoRam_00_9(),
  function ActionValue#(Struct19) getRs_infoRam_00_8(),
  function ActionValue#(Struct19) getRs_infoRam_00_7(),
  function ActionValue#(Struct19) getRs_infoRam_00_6(),
  function ActionValue#(Struct19) getRs_infoRam_00_5(),
  function ActionValue#(Struct19) getRs_infoRam_00_4(),
  function ActionValue#(Struct19) getRs_infoRam_00_3(),
  function ActionValue#(Struct19) getRs_infoRam_00_2(),
  function ActionValue#(Struct19) getRs_infoRam_00_1(),
  function ActionValue#(Struct19) getRs_infoRam_00_0()) (Module133);
    Reg#(Bit#(2)) readStage_00 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_00 <- mkReg(unpack(0));
    Reg#(Struct3) readLine_00 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_00 <- mkReg(unpack(0));
    Reg#(Struct3) writeLine_00 <- mkReg(unpack(0));
    Reg#(Vector#(8, Struct18)) victims_00 <- mkReg(unpack(0));
    Reg#(Struct3) victimLine_00 <- mkReg(unpack(0));
    Reg#(Bit#(4)) victimWay_00 <- mkReg(unpack(0));

    rule read_tagmatch_00;
        let x_0 = (readStage_00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_00);
        Bit#(51) x_2 = ((x_1)[63:13]);
        Bit#(10) x_3 = ((x_1)[12:3]);
        Vector#(16, Struct19) x_4 =
        ((Vector#(16, Struct19))'(vec(Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_00_0();
        Vector#(16, Struct19) x_6 = (update (x_4, (Bit#(4))'(4'h0), x_5));
        let x_7 <- getRs_infoRam_00_1();
        Vector#(16, Struct19) x_8 = (update (x_6, (Bit#(4))'(4'h1), x_7));
        let x_9 <- getRs_infoRam_00_2();
        Vector#(16, Struct19) x_10 = (update (x_8, (Bit#(4))'(4'h2), x_9));

        let x_11 <- getRs_infoRam_00_3();
        Vector#(16, Struct19) x_12 = (update (x_10, (Bit#(4))'(4'h3), x_11));

        let x_13 <- getRs_infoRam_00_4();
        Vector#(16, Struct19) x_14 = (update (x_12, (Bit#(4))'(4'h4), x_13));

        let x_15 <- getRs_infoRam_00_5();
        Vector#(16, Struct19) x_16 = (update (x_14, (Bit#(4))'(4'h5), x_15));

        let x_17 <- getRs_infoRam_00_6();
        Vector#(16, Struct19) x_18 = (update (x_16, (Bit#(4))'(4'h6), x_17));

        let x_19 <- getRs_infoRam_00_7();
        Vector#(16, Struct19) x_20 = (update (x_18, (Bit#(4))'(4'h7), x_19));

        let x_21 <- getRs_infoRam_00_8();
        Vector#(16, Struct19) x_22 = (update (x_20, (Bit#(4))'(4'h8), x_21));

        let x_23 <- getRs_infoRam_00_9();
        Vector#(16, Struct19) x_24 = (update (x_22, (Bit#(4))'(4'h9), x_23));

        let x_25 <- getRs_infoRam_00_10();
        Vector#(16, Struct19) x_26 = (update (x_24, (Bit#(4))'(4'ha), x_25));

        let x_27 <- getRs_infoRam_00_11();
        Vector#(16, Struct19) x_28 = (update (x_26, (Bit#(4))'(4'hb), x_27));

        let x_29 <- getRs_infoRam_00_12();
        Vector#(16, Struct19) x_30 = (update (x_28, (Bit#(4))'(4'hc), x_29));

        let x_31 <- getRs_infoRam_00_13();
        Vector#(16, Struct19) x_32 = (update (x_30, (Bit#(4))'(4'hd), x_31));

        let x_33 <- getRs_infoRam_00_14();
        Vector#(16, Struct19) x_34 = (update (x_32, (Bit#(4))'(4'he), x_33));

        let x_35 <- getRs_infoRam_00_15();
        Vector#(16, Struct19) x_36 = (update (x_34, (Bit#(4))'(4'hf), x_35));

        Struct20 x_37 = (((((x_36)[(Bit#(4))'(4'h0)]).tag) == (x_2) ?
        (Struct20 {tm_hit : (Bool)'(True), tm_way : (Bit#(4))'(4'h0),
        tm_value : ((x_36)[(Bit#(4))'(4'h0)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h1)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h1), tm_value :
        ((x_36)[(Bit#(4))'(4'h1)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h2)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h2), tm_value :
        ((x_36)[(Bit#(4))'(4'h2)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h3)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h3), tm_value :
        ((x_36)[(Bit#(4))'(4'h3)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h4)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h4), tm_value :
        ((x_36)[(Bit#(4))'(4'h4)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h5)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h5), tm_value :
        ((x_36)[(Bit#(4))'(4'h5)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h6)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h6), tm_value :
        ((x_36)[(Bit#(4))'(4'h6)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h7)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h7), tm_value :
        ((x_36)[(Bit#(4))'(4'h7)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h8)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h8), tm_value :
        ((x_36)[(Bit#(4))'(4'h8)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h9)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h9), tm_value :
        ((x_36)[(Bit#(4))'(4'h9)]).value}) :
        (((((x_36)[(Bit#(4))'(4'ha)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'ha), tm_value :
        ((x_36)[(Bit#(4))'(4'ha)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hb)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hb), tm_value :
        ((x_36)[(Bit#(4))'(4'hb)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hc)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hc), tm_value :
        ((x_36)[(Bit#(4))'(4'hc)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hd)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hd), tm_value :
        ((x_36)[(Bit#(4))'(4'hd)]).value}) :
        (((((x_36)[(Bit#(4))'(4'he)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'he), tm_value :
        ((x_36)[(Bit#(4))'(4'he)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hf)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hf), tm_value :
        ((x_36)[(Bit#(4))'(4'hf)]).value}) :
        ((Struct20)'(Struct20 {tm_hit: False, tm_way: 4'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))))))))))))))))))))))))))));

        readLine_00 <= Struct3 {addr : x_1, info_hit : (x_37).tm_hit,
        info_way : (x_37).tm_way, info_write : (Bool)'(False), info :
        (x_37).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_37).tm_hit) begin

            readStage_00 <= (Bit#(2))'(2'h2);
            let x_38 <- putRq_dataRam_00(Struct21 {write : (Bool)'(False),
            addr : {(x_3),((x_37).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_00 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_00;
        let x_0 = (readStage_00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_00 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_00();
        let x_2 = (readLine_00);
        readLine_00 <= Struct3 {addr : (x_2).addr, info_hit : (x_2).info_hit,
        info_way : (x_2).info_way, info_write : (x_2).info_write, info :
        (x_2).info, value_write : (Bool)'(False), value : x_1};

    endrule

    rule write_info_hit_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_00);
        when ((x_1).info_hit, noAction);
        writeStage_00 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(10) x_4 = ((x_2)[12:3]);
        Bit#(4) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct22 x_6 = (Struct22 {write : (Bool)'(True), addr : x_4,
            datain : Struct19 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(4))'(4'h0))) begin
            let x_7 <- putRq_infoRam_00_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h1))) begin
            let x_9 <- putRq_infoRam_00_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h2))) begin
            let x_11 <- putRq_infoRam_00_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h3))) begin
            let x_13 <- putRq_infoRam_00_3(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h4))) begin
            let x_15 <- putRq_infoRam_00_4(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h5))) begin
            let x_17 <- putRq_infoRam_00_5(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h6))) begin
            let x_19 <- putRq_infoRam_00_6(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h7))) begin
            let x_21 <- putRq_infoRam_00_7(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h8))) begin
            let x_23 <- putRq_infoRam_00_8(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h9))) begin
            let x_25 <- putRq_infoRam_00_9(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'ha))) begin
            let x_27 <- putRq_infoRam_00_10(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hb))) begin
            let x_29 <- putRq_infoRam_00_11(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hc))) begin
            let x_31 <- putRq_infoRam_00_12(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hd))) begin
            let x_33 <- putRq_infoRam_00_13(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'he))) begin
            let x_35 <- putRq_infoRam_00_14(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hf))) begin
            let x_37 <- putRq_infoRam_00_15(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_40 <- putRq_dataRam_00(Struct21 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_00);
        when (! ((x_1).info_hit), noAction);
        writeStage_00 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(10) x_3 = ((x_2)[12:3]);
        Struct22 x_4 = (Struct22 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct19)'(Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_00_0(x_4);
        let x_6 <- putRq_infoRam_00_1(x_4);
        let x_7 <- putRq_infoRam_00_2(x_4);
        let x_8 <- putRq_infoRam_00_3(x_4);
        let x_9 <- putRq_infoRam_00_4(x_4);
        let x_10 <- putRq_infoRam_00_5(x_4);
        let x_11 <- putRq_infoRam_00_6(x_4);
        let x_12 <- putRq_infoRam_00_7(x_4);
        let x_13 <- putRq_infoRam_00_8(x_4);
        let x_14 <- putRq_infoRam_00_9(x_4);
        let x_15 <- putRq_infoRam_00_10(x_4);
        let x_16 <- putRq_infoRam_00_11(x_4);
        let x_17 <- putRq_infoRam_00_12(x_4);
        let x_18 <- putRq_infoRam_00_13(x_4);
        let x_19 <- putRq_infoRam_00_14(x_4);
        let x_20 <- putRq_infoRam_00_15(x_4);

    endrule

    rule write_info_miss_rep_rs_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_00 <= (Bit#(3))'(3'h3);
        Vector#(16, Struct19) x_1 =
        ((Vector#(16, Struct19))'(vec(Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_00_0();
        Vector#(16, Struct19) x_3 = (update (x_1, (Bit#(4))'(4'h0), x_2));
        let x_4 <- getRs_infoRam_00_1();
        Vector#(16, Struct19) x_5 = (update (x_3, (Bit#(4))'(4'h1), x_4));
        let x_6 <- getRs_infoRam_00_2();
        Vector#(16, Struct19) x_7 = (update (x_5, (Bit#(4))'(4'h2), x_6));
        let x_8 <- getRs_infoRam_00_3();
        Vector#(16, Struct19) x_9 = (update (x_7, (Bit#(4))'(4'h3), x_8));
        let x_10 <- getRs_infoRam_00_4();
        Vector#(16, Struct19) x_11 = (update (x_9, (Bit#(4))'(4'h4), x_10));

        let x_12 <- getRs_infoRam_00_5();
        Vector#(16, Struct19) x_13 = (update (x_11, (Bit#(4))'(4'h5), x_12));

        let x_14 <- getRs_infoRam_00_6();
        Vector#(16, Struct19) x_15 = (update (x_13, (Bit#(4))'(4'h6), x_14));

        let x_16 <- getRs_infoRam_00_7();
        Vector#(16, Struct19) x_17 = (update (x_15, (Bit#(4))'(4'h7), x_16));

        let x_18 <- getRs_infoRam_00_8();
        Vector#(16, Struct19) x_19 = (update (x_17, (Bit#(4))'(4'h8), x_18));

        let x_20 <- getRs_infoRam_00_9();
        Vector#(16, Struct19) x_21 = (update (x_19, (Bit#(4))'(4'h9), x_20));

        let x_22 <- getRs_infoRam_00_10();
        Vector#(16, Struct19) x_23 = (update (x_21, (Bit#(4))'(4'ha), x_22));

        let x_24 <- getRs_infoRam_00_11();
        Vector#(16, Struct19) x_25 = (update (x_23, (Bit#(4))'(4'hb), x_24));

        let x_26 <- getRs_infoRam_00_12();
        Vector#(16, Struct19) x_27 = (update (x_25, (Bit#(4))'(4'hc), x_26));

        let x_28 <- getRs_infoRam_00_13();
        Vector#(16, Struct19) x_29 = (update (x_27, (Bit#(4))'(4'hd), x_28));

        let x_30 <- getRs_infoRam_00_14();
        Vector#(16, Struct19) x_31 = (update (x_29, (Bit#(4))'(4'he), x_30));

        let x_32 <- getRs_infoRam_00_15();
        Vector#(16, Struct19) x_33 = (update (x_31, (Bit#(4))'(4'hf), x_32));

        Bit#(4) x_34 = ((((((x_33)[(Bit#(4))'(4'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h0)) :
        ((((((x_33)[(Bit#(4))'(4'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h1)) :
        ((((((x_33)[(Bit#(4))'(4'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h2)) :
        ((((((x_33)[(Bit#(4))'(4'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h3)) :
        ((((((x_33)[(Bit#(4))'(4'h4)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h4)) :
        ((((((x_33)[(Bit#(4))'(4'h5)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h5)) :
        ((((((x_33)[(Bit#(4))'(4'h6)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h6)) :
        ((((((x_33)[(Bit#(4))'(4'h7)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h7)) :
        ((((((x_33)[(Bit#(4))'(4'h8)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h8)) :
        ((((((x_33)[(Bit#(4))'(4'h9)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h9)) :
        ((((((x_33)[(Bit#(4))'(4'ha)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'ha)) :
        ((((((x_33)[(Bit#(4))'(4'hb)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hb)) :
        ((((((x_33)[(Bit#(4))'(4'hc)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hc)) :
        ((((((x_33)[(Bit#(4))'(4'hd)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hd)) :
        ((((((x_33)[(Bit#(4))'(4'he)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'he)) :
        ((((((x_33)[(Bit#(4))'(4'hf)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hf)) :
        ((Bit#(4))'(4'h0))))))))))))))))))))))))))))))))));
        let x_35 = (writeLine_00);
        Bit#(64) x_36 = ((x_35).addr);
        Bit#(10) x_37 = ((x_36)[12:3]);
        Struct19 x_38 = ((x_33)[x_34]);
        Bit#(51) x_39 = ((x_38).tag);
        Struct4 x_40 = ((x_38).value);
        victimWay_00 <= x_34;
        victimLine_00 <= Struct3 {addr :
        {(x_39),({(x_37),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(4))'(4'h0), info_write : (Bool)'(False), info :
        x_40, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_41 <- putRq_dataRam_00(Struct21 {write : (Bool)'(False), addr :
        {(x_37),(x_34)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_00);
        writeStage_00 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(10) x_4 = ((x_2)[12:3]);
        let x_5 = (victimWay_00);
        let x_6 = (victims_00);
        when ((! (((x_6)[(Bit#(3))'(3'h7)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h6)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h5)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h4)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(3))'(3'h0)]).victim_valid)))))))), noAction);
        Bit#(3) x_7 = ((((x_6)[(Bit#(3))'(3'h7)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h6)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h5)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h4)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h3)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h2)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h1)]).victim_valid ? ((Bit#(3))'(3'h0)) :
        ((Bit#(3))'(3'h1)))) : ((Bit#(3))'(3'h2)))) : ((Bit#(3))'(3'h3)))) :
        ((Bit#(3))'(3'h4)))) : ((Bit#(3))'(3'h5)))) : ((Bit#(3))'(3'h6)))) :
        ((Bit#(3))'(3'h7))));
        let x_8 <- getRs_dataRam_00();
        let x_9 = (victimLine_00);
        victims_00 <= update (x_6, x_7, Struct18 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct3 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_00 <= Struct3 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct22 x_10 = (Struct22 {write : (Bool)'(True), addr : x_4,
            datain : Struct19 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(4))'(4'h0))) begin
            let x_11 <- putRq_infoRam_00_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h1))) begin
            let x_13 <- putRq_infoRam_00_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h2))) begin
            let x_15 <- putRq_infoRam_00_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h3))) begin
            let x_17 <- putRq_infoRam_00_3(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h4))) begin
            let x_19 <- putRq_infoRam_00_4(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h5))) begin
            let x_21 <- putRq_infoRam_00_5(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h6))) begin
            let x_23 <- putRq_infoRam_00_6(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h7))) begin
            let x_25 <- putRq_infoRam_00_7(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h8))) begin
            let x_27 <- putRq_infoRam_00_8(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h9))) begin
            let x_29 <- putRq_infoRam_00_9(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'ha))) begin
            let x_31 <- putRq_infoRam_00_10(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hb))) begin
            let x_33 <- putRq_infoRam_00_11(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hc))) begin
            let x_35 <- putRq_infoRam_00_12(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hd))) begin
            let x_37 <- putRq_infoRam_00_13(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'he))) begin
            let x_39 <- putRq_infoRam_00_14(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hf))) begin
            let x_41 <- putRq_infoRam_00_15(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_44 <- putRq_dataRam_00(Struct21 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_00_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_00);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_00);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_00);
        Struct18 x_4 = ((x_3)[(Bit#(3))'(3'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_00 <= (Bit#(2))'(2'h3);
        readLine_00 <= (x_4).victim_line;

        end else begin

            Struct18 x_5 = ((x_3)[(Bit#(3))'(3'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_00 <= (Bit#(2))'(2'h3);
                readLine_00 <= (x_5).victim_line;

            end else begin

                Struct18 x_6 = ((x_3)[(Bit#(3))'(3'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_00 <= (Bit#(2))'(2'h3);
                    readLine_00 <= (x_6).victim_line;

                end else begin

                    Struct18 x_7 = ((x_3)[(Bit#(3))'(3'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_00 <= (Bit#(2))'(2'h3);
                        readLine_00 <= (x_7).victim_line;

                    end else begin

                        Struct18 x_8 = ((x_3)[(Bit#(3))'(3'h4)]);
                        if (((x_8).victim_valid) &&
                        ((((x_8).victim_line).addr) == (x_0))) begin

                            readStage_00 <= (Bit#(2))'(2'h3);
                            readLine_00 <= (x_8).victim_line;

                        end else begin

                            Struct18 x_9 = ((x_3)[(Bit#(3))'(3'h5)]);
                            if (((x_9).victim_valid) &&
                            ((((x_9).victim_line).addr) == (x_0))) begin

                                readStage_00 <= (Bit#(2))'(2'h3);
                                readLine_00 <= (x_9).victim_line;

                            end else begin

                                Struct18 x_10 = ((x_3)[(Bit#(3))'(3'h6)]);
                                if (((x_10).victim_valid) &&
                                ((((x_10).victim_line).addr) == (x_0))) begin

                                    readStage_00 <= (Bit#(2))'(2'h3);

                                    readLine_00 <= (x_10).victim_line;

                                end else begin

                                    Struct18 x_11 = ((x_3)[(Bit#(3))'(3'h7)]);

                                    if (((x_11).victim_valid) &&
                                    ((((x_11).victim_line).addr) == (x_0)))
                                    begin

                                        readStage_00 <= (Bit#(2))'(2'h3);

                                        readLine_00 <= (x_11).victim_line;

                                    end else begin

                                        readStage_00 <= (Bit#(2))'(2'h1);

                                        readAddr_00 <= x_0;
                                        Bit#(10) x_12 = ((x_0)[12:3]);

                                        Struct22 x_13 = (Struct22 {write :
                                        (Bool)'(False), addr : x_12, datain :
                                        (Struct19)'(Struct19 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                                        let x_14 <- putRq_infoRam_00_0(x_13);

                                        let x_15 <- putRq_infoRam_00_1(x_13);

                                        let x_16 <- putRq_infoRam_00_2(x_13);

                                        let x_17 <- putRq_infoRam_00_3(x_13);

                                        let x_18 <- putRq_infoRam_00_4(x_13);

                                        let x_19 <- putRq_infoRam_00_5(x_13);

                                        let x_20 <- putRq_infoRam_00_6(x_13);

                                        let x_21 <- putRq_infoRam_00_7(x_13);

                                        let x_22 <- putRq_infoRam_00_8(x_13);

                                        let x_23 <- putRq_infoRam_00_9(x_13);

                                        let x_24 <-
                                        putRq_infoRam_00_10(x_13);
                                        let x_25 <-
                                        putRq_infoRam_00_11(x_13);
                                        let x_26 <-
                                        putRq_infoRam_00_12(x_13);
                                        let x_27 <-
                                        putRq_infoRam_00_13(x_13);
                                        let x_28 <-
                                        putRq_infoRam_00_14(x_13);
                                        let x_29 <-
                                        putRq_infoRam_00_15(x_13);

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct3) cache_00_readRs ();
        let x_1 = (readStage_00);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_00 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_00);
        return x_2;
    endmethod

    method Action cache_00_writeRq (Struct3 x_0);
        let x_1 = (readStage_00);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_00);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_00);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct18 x_5 = ((x_3)[(Bit#(3))'(3'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct3 x_6 = (Struct3 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h1)));

            writeLine_00 <= x_6;
            victims_00 <= update (x_3, (Bit#(3))'(3'h0), Struct18
            {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h0), victim_line :
            x_6});

        end else begin

            Struct18 x_7 = ((x_3)[(Bit#(3))'(3'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct3 x_8 = (Struct3 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_00 <= x_8;
                victims_00 <= update (x_3, (Bit#(3))'(3'h1), Struct18
                {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h1),
                victim_line : x_8});

            end else begin

                Struct18 x_9 = ((x_3)[(Bit#(3))'(3'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct3 x_10 = (Struct3 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_00 <= x_10;
                    victims_00 <= update (x_3, (Bit#(3))'(3'h2), Struct18
                    {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h2),
                    victim_line : x_10});

                end else begin

                    Struct18 x_11 = ((x_3)[(Bit#(3))'(3'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct3 x_12 = (Struct3 {addr : (x_0).addr, info_hit
                        : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_00 <= x_12;
                        victims_00 <= update (x_3, (Bit#(3))'(3'h3), Struct18
                        {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h3),
                        victim_line : x_12});

                    end else begin

                        Struct18 x_13 = ((x_3)[(Bit#(3))'(3'h4)]);
                        if (((x_13).victim_valid) &&
                        ((((x_13).victim_line).addr) == ((x_0).addr))) begin

                            Struct3 x_14 = (Struct3 {addr : (x_0).addr,
                            info_hit : (Bool)'(False), info_way :
                            (x_0).info_way, info_write : (x_0).info_write,
                            info : (x_0).info, value_write :
                            (x_0).value_write, value : (x_0).value});

                            writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                            ((Bit#(3))'(3'h1)));
                            writeLine_00 <= x_14;
                            victims_00 <= update (x_3, (Bit#(3))'(3'h4),
                            Struct18 {victim_valid : x_4, victim_idx :
                            (Bit#(3))'(3'h4), victim_line : x_14});

                        end else begin

                            Struct18 x_15 = ((x_3)[(Bit#(3))'(3'h5)]);
                            if (((x_15).victim_valid) &&
                            ((((x_15).victim_line).addr) == ((x_0).addr)))
                            begin

                                Struct3 x_16 = (Struct3 {addr : (x_0).addr,
                                info_hit : (Bool)'(False), info_way :
                                (x_0).info_way, info_write :
                                (x_0).info_write, info : (x_0).info,
                                value_write : (x_0).value_write, value :
                                (x_0).value});
                                writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                                ((Bit#(3))'(3'h1)));
                                writeLine_00 <= x_16;
                                victims_00 <= update (x_3, (Bit#(3))'(3'h5),
                                Struct18 {victim_valid : x_4, victim_idx :
                                (Bit#(3))'(3'h5), victim_line : x_16});

                            end else begin

                                Struct18 x_17 = ((x_3)[(Bit#(3))'(3'h6)]);
                                if (((x_17).victim_valid) &&
                                ((((x_17).victim_line).addr) ==
                                ((x_0).addr))) begin

                                    Struct3 x_18 = (Struct3 {addr :
                                    (x_0).addr, info_hit : (Bool)'(False),
                                    info_way : (x_0).info_way, info_write :
                                    (x_0).info_write, info : (x_0).info,
                                    value_write : (x_0).value_write, value :
                                    (x_0).value});
                                    writeStage_00 <= (x_4 ?
                                    ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h1)));

                                    writeLine_00 <= x_18;
                                    victims_00 <= update (x_3,
                                    (Bit#(3))'(3'h6), Struct18 {victim_valid
                                    : x_4, victim_idx : (Bit#(3))'(3'h6),
                                    victim_line : x_18});

                                end else begin

                                    Struct18 x_19 = ((x_3)[(Bit#(3))'(3'h7)]);

                                    if (((x_19).victim_valid) &&
                                    ((((x_19).victim_line).addr) ==
                                    ((x_0).addr))) begin

                                        Struct3 x_20 = (Struct3 {addr :
                                        (x_0).addr, info_hit :
                                        (Bool)'(False), info_way :
                                        (x_0).info_way, info_write :
                                        (x_0).info_write, info : (x_0).info,
                                        value_write : (x_0).value_write,
                                        value : (x_0).value});
                                        writeStage_00 <= (x_4 ?
                                        ((Bit#(3))'(3'h7)) :
                                        ((Bit#(3))'(3'h1)));
                                        writeLine_00 <= x_20;
                                        victims_00 <= update (x_3,
                                        (Bit#(3))'(3'h7), Struct18
                                        {victim_valid : x_4, victim_idx :
                                        (Bit#(3))'(3'h7), victim_line :
                                        x_20});

                                    end else begin

                                        writeStage_00 <= (Bit#(3))'(3'h1);

                                        writeLine_00 <= x_0;

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct3) cache_00_writeRs ();
        let x_1 = (writeStage_00);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_00 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_00);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_00_hasVictimSlot ();
        let x_1 = (victims_00);
        Bool x_2 = ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) ||
        (((x_1)[(Bit#(3))'(3'h0)]).victim_valid))))))));
        return x_2;
    endmethod

    method ActionValue#(Struct3) cache_00_getVictim ();
        let x_1 = (victims_00);
        when ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) ||
        (((x_1)[(Bit#(3))'(3'h0)]).victim_valid))))))), noAction);
        Struct3 x_2 = ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h7)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h6)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h5)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h4)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h3)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h2)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h1)]).victim_line) :
        (((x_1)[(Bit#(3))'(3'h0)]).victim_line)))))))))))))));
        return x_2;
    endmethod

    method Action cache_00_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_00);
        Struct18 x_2 = ((x_1)[(Bit#(3))'(3'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_00 <= update (x_1, (Bit#(3))'(3'h0),
            (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct18 x_3 = ((x_1)[(Bit#(3))'(3'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_00 <= update (x_1, (Bit#(3))'(3'h1),
                (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct18 x_4 = ((x_1)[(Bit#(3))'(3'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_00 <= update (x_1, (Bit#(3))'(3'h2),
                    (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct18 x_5 = ((x_1)[(Bit#(3))'(3'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_00 <= update (x_1, (Bit#(3))'(3'h3),
                        (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                        Struct18 x_6 = ((x_1)[(Bit#(3))'(3'h4)]);
                        if (((x_6).victim_valid) &&
                        ((((x_6).victim_line).addr) == (x_0))) begin

                            victims_00 <= update (x_1, (Bit#(3))'(3'h4),
                            (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                        end else begin

                            Struct18 x_7 = ((x_1)[(Bit#(3))'(3'h5)]);
                            if (((x_7).victim_valid) &&
                            ((((x_7).victim_line).addr) == (x_0))) begin

                                victims_00 <= update (x_1, (Bit#(3))'(3'h5),
                                (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                            end else begin

                                Struct18 x_8 = ((x_1)[(Bit#(3))'(3'h6)]);
                                if (((x_8).victim_valid) &&
                                ((((x_8).victim_line).addr) == (x_0))) begin

                                    victims_00 <= update (x_1,
                                    (Bit#(3))'(3'h6),
                                    (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                                end else begin

                                    Struct18 x_9 = ((x_1)[(Bit#(3))'(3'h7)]);

                                    if (((x_9).victim_valid) &&
                                    ((((x_9).victim_line).addr) == (x_0)))
                                    begin

                                        victims_00 <= update (x_1,
                                        (Bit#(3))'(3'h7),
                                        (Struct18)'(Struct18 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                                    end else begin

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

endmodule

interface Module134;
    method Action makeEnq_parentChildren00 (Struct10 x_0);
    method Action broadcast_parentChildren00 (Struct13 x_0);

endinterface


module mkModule134#(function Action enq_fifo0002(Struct2 _),
  function Action enq_fifo0012(Struct2 _),
  function Action enq_fifo0022(Struct2 _),
  function Action enq_fifo0032(Struct2 _),
  function Action enq_fifo001(Struct2 _),
  function Action enq_fifo000(Struct2 _)) (Module134);

    // No rules in this module

    method Action makeEnq_parentChildren00 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo000((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo001((x_0).enq_msg);

            end else begin

                Bit#(2) x_3 = ((x_0).enq_ch_idx);
                Struct2 x_4 = ((x_0).enq_msg);
                if ((x_3) == ((Bit#(2))'(2'h3))) begin
                let x_5 <- enq_fifo0032(x_4);

                end else begin

                    if ((x_3) == ((Bit#(2))'(2'h2))) begin
                    let x_6 <- enq_fifo0022(x_4);

                    end else begin

                        if ((x_3) == ((Bit#(2))'(2'h1))) begin
                        let x_7 <- enq_fifo0012(x_4);

                        end else begin

                            if ((x_3) == ((Bit#(2))'(2'h0))) begin
                            let x_8 <- enq_fifo0002(x_4);

                            end else begin

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method Action broadcast_parentChildren00 (Struct13 x_0);
        Bit#(4) x_1 = ((x_0).cs_inds);
        Struct2 x_2 = ((x_0).cs_msg);
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == (x_1))
        begin
        let x_3 <- enq_fifo0032(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == (x_1))
        begin
        let x_5 <- enq_fifo0022(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == (x_1))
        begin
        let x_7 <- enq_fifo0012(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == (x_1))
        begin
        let x_9 <- enq_fifo0002(x_2);

        end else begin

        end

    endmethod

endmodule

interface Module135;
    method Action cache_000_readRq (Bit#(64) x_0);
    method ActionValue#(Struct24) cache_000_readRs ();
    method Action cache_000_writeRq (Struct24 x_0);
    method ActionValue#(Struct24) cache_000_writeRs ();
    method ActionValue#(Bool) cache_000_hasVictimSlot ();
    method ActionValue#(Struct24) cache_000_getVictim ();
    method Action cache_000_removeVictim (Bit#(64) x_0);

endinterface


module mkModule135#(function Action putRq_infoRam_000_7(Struct29 _),
  function Action putRq_infoRam_000_6(Struct29 _),
  function Action putRq_infoRam_000_5(Struct29 _),
  function Action putRq_infoRam_000_4(Struct29 _),
  function Action putRq_infoRam_000_3(Struct29 _),
  function Action putRq_infoRam_000_2(Struct29 _),
  function Action putRq_infoRam_000_1(Struct29 _),
  function Action putRq_infoRam_000_0(Struct29 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_000(),
  function Action putRq_dataRam_000(Struct28 _),
  function ActionValue#(Struct26) getRs_infoRam_000_7(),
  function ActionValue#(Struct26) getRs_infoRam_000_6(),
  function ActionValue#(Struct26) getRs_infoRam_000_5(),
  function ActionValue#(Struct26) getRs_infoRam_000_4(),
  function ActionValue#(Struct26) getRs_infoRam_000_3(),
  function ActionValue#(Struct26) getRs_infoRam_000_2(),
  function ActionValue#(Struct26) getRs_infoRam_000_1(),
  function ActionValue#(Struct26) getRs_infoRam_000_0()) (Module135);
    Reg#(Bit#(2)) readStage_000 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_000 <- mkReg(unpack(0));
    Reg#(Struct24) readLine_000 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_000 <- mkReg(unpack(0));
    Reg#(Struct24) writeLine_000 <- mkReg(unpack(0));
    Reg#(Vector#(8, Struct25)) victims_000 <- mkReg(unpack(0));
    Reg#(Struct24) victimLine_000 <- mkReg(unpack(0));
    Reg#(Bit#(3)) victimWay_000 <- mkReg(unpack(0));

    rule read_tagmatch_000;
        let x_0 = (readStage_000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_000);
        Bit#(53) x_2 = ((x_1)[63:11]);
        Bit#(8) x_3 = ((x_1)[10:3]);
        Vector#(8, Struct26) x_4 =
        ((Vector#(8, Struct26))'(vec(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_000_0();
        Vector#(8, Struct26) x_6 = (update (x_4, (Bit#(3))'(3'h0), x_5));
        let x_7 <- getRs_infoRam_000_1();
        Vector#(8, Struct26) x_8 = (update (x_6, (Bit#(3))'(3'h1), x_7));
        let x_9 <- getRs_infoRam_000_2();
        Vector#(8, Struct26) x_10 = (update (x_8, (Bit#(3))'(3'h2), x_9));
        let x_11 <- getRs_infoRam_000_3();
        Vector#(8, Struct26) x_12 = (update (x_10, (Bit#(3))'(3'h3), x_11));

        let x_13 <- getRs_infoRam_000_4();
        Vector#(8, Struct26) x_14 = (update (x_12, (Bit#(3))'(3'h4), x_13));

        let x_15 <- getRs_infoRam_000_5();
        Vector#(8, Struct26) x_16 = (update (x_14, (Bit#(3))'(3'h5), x_15));

        let x_17 <- getRs_infoRam_000_6();
        Vector#(8, Struct26) x_18 = (update (x_16, (Bit#(3))'(3'h6), x_17));

        let x_19 <- getRs_infoRam_000_7();
        Vector#(8, Struct26) x_20 = (update (x_18, (Bit#(3))'(3'h7), x_19));

        Struct27 x_21 = (((((x_20)[(Bit#(3))'(3'h0)]).tag) == (x_2) ?
        (Struct27 {tm_hit : (Bool)'(True), tm_way : (Bit#(3))'(3'h0),
        tm_value : ((x_20)[(Bit#(3))'(3'h0)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h1)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h1), tm_value :
        ((x_20)[(Bit#(3))'(3'h1)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h2)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h2), tm_value :
        ((x_20)[(Bit#(3))'(3'h2)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h3)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h3), tm_value :
        ((x_20)[(Bit#(3))'(3'h3)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h4)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h4), tm_value :
        ((x_20)[(Bit#(3))'(3'h4)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h5)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h5), tm_value :
        ((x_20)[(Bit#(3))'(3'h5)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h6)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h6), tm_value :
        ((x_20)[(Bit#(3))'(3'h6)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h7)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h7), tm_value :
        ((x_20)[(Bit#(3))'(3'h7)]).value}) :
        ((Struct27)'(Struct27 {tm_hit: False, tm_way: 3'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))))))))))));

        readLine_000 <= Struct24 {addr : x_1, info_hit : (x_21).tm_hit,
        info_way : (x_21).tm_way, info_write : (Bool)'(False), info :
        (x_21).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_21).tm_hit) begin

            readStage_000 <= (Bit#(2))'(2'h2);
            let x_22 <- putRq_dataRam_000(Struct28 {write : (Bool)'(False),
            addr : {(x_3),((x_21).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_000 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_000;
        let x_0 = (readStage_000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_000 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_000();
        let x_2 = (readLine_000);
        readLine_000 <= Struct24 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_000);
        when ((x_1).info_hit, noAction);
        writeStage_000 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(53) x_3 = ((x_2)[63:11]);
        Bit#(8) x_4 = ((x_2)[10:3]);
        Bit#(3) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct29 x_6 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(3))'(3'h0))) begin
            let x_7 <- putRq_infoRam_000_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h1))) begin
            let x_9 <- putRq_infoRam_000_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h2))) begin
            let x_11 <- putRq_infoRam_000_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h3))) begin
            let x_13 <- putRq_infoRam_000_3(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h4))) begin
            let x_15 <- putRq_infoRam_000_4(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h5))) begin
            let x_17 <- putRq_infoRam_000_5(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h6))) begin
            let x_19 <- putRq_infoRam_000_6(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h7))) begin
            let x_21 <- putRq_infoRam_000_7(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_24 <- putRq_dataRam_000(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_000);
        when (! ((x_1).info_hit), noAction);
        writeStage_000 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(8) x_3 = ((x_2)[10:3]);
        Struct29 x_4 = (Struct29 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct26)'(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_000_0(x_4);
        let x_6 <- putRq_infoRam_000_1(x_4);
        let x_7 <- putRq_infoRam_000_2(x_4);
        let x_8 <- putRq_infoRam_000_3(x_4);
        let x_9 <- putRq_infoRam_000_4(x_4);
        let x_10 <- putRq_infoRam_000_5(x_4);
        let x_11 <- putRq_infoRam_000_6(x_4);
        let x_12 <- putRq_infoRam_000_7(x_4);

    endrule

    rule write_info_miss_rep_rs_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_000 <= (Bit#(3))'(3'h3);
        Vector#(8, Struct26) x_1 =
        ((Vector#(8, Struct26))'(vec(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_000_0();
        Vector#(8, Struct26) x_3 = (update (x_1, (Bit#(3))'(3'h0), x_2));
        let x_4 <- getRs_infoRam_000_1();
        Vector#(8, Struct26) x_5 = (update (x_3, (Bit#(3))'(3'h1), x_4));
        let x_6 <- getRs_infoRam_000_2();
        Vector#(8, Struct26) x_7 = (update (x_5, (Bit#(3))'(3'h2), x_6));
        let x_8 <- getRs_infoRam_000_3();
        Vector#(8, Struct26) x_9 = (update (x_7, (Bit#(3))'(3'h3), x_8));
        let x_10 <- getRs_infoRam_000_4();
        Vector#(8, Struct26) x_11 = (update (x_9, (Bit#(3))'(3'h4), x_10));

        let x_12 <- getRs_infoRam_000_5();
        Vector#(8, Struct26) x_13 = (update (x_11, (Bit#(3))'(3'h5), x_12));

        let x_14 <- getRs_infoRam_000_6();
        Vector#(8, Struct26) x_15 = (update (x_13, (Bit#(3))'(3'h6), x_14));

        let x_16 <- getRs_infoRam_000_7();
        Vector#(8, Struct26) x_17 = (update (x_15, (Bit#(3))'(3'h7), x_16));

        Bit#(3) x_18 = ((((((x_17)[(Bit#(3))'(3'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h0)) :
        ((((((x_17)[(Bit#(3))'(3'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h1)) :
        ((((((x_17)[(Bit#(3))'(3'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h2)) :
        ((((((x_17)[(Bit#(3))'(3'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h3)) :
        ((((((x_17)[(Bit#(3))'(3'h4)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h4)) :
        ((((((x_17)[(Bit#(3))'(3'h5)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h5)) :
        ((((((x_17)[(Bit#(3))'(3'h6)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h6)) :
        ((((((x_17)[(Bit#(3))'(3'h7)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h7)) :
        ((Bit#(3))'(3'h0))))))))))))))))));
        let x_19 = (writeLine_000);
        Bit#(64) x_20 = ((x_19).addr);
        Bit#(8) x_21 = ((x_20)[10:3]);
        Struct26 x_22 = ((x_17)[x_18]);
        Bit#(53) x_23 = ((x_22).tag);
        Struct4 x_24 = ((x_22).value);
        victimWay_000 <= x_18;
        victimLine_000 <= Struct24 {addr :
        {(x_23),({(x_21),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(3))'(3'h0), info_write : (Bool)'(False), info :
        x_24, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_25 <- putRq_dataRam_000(Struct28 {write : (Bool)'(False), addr
        : {(x_21),(x_18)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_000);
        writeStage_000 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(53) x_3 = ((x_2)[63:11]);
        Bit#(8) x_4 = ((x_2)[10:3]);
        let x_5 = (victimWay_000);
        let x_6 = (victims_000);
        when ((! (((x_6)[(Bit#(3))'(3'h7)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h6)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h5)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h4)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(3))'(3'h0)]).victim_valid)))))))), noAction);
        Bit#(3) x_7 = ((((x_6)[(Bit#(3))'(3'h7)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h6)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h5)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h4)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h3)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h2)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h1)]).victim_valid ? ((Bit#(3))'(3'h0)) :
        ((Bit#(3))'(3'h1)))) : ((Bit#(3))'(3'h2)))) : ((Bit#(3))'(3'h3)))) :
        ((Bit#(3))'(3'h4)))) : ((Bit#(3))'(3'h5)))) : ((Bit#(3))'(3'h6)))) :
        ((Bit#(3))'(3'h7))));
        let x_8 <- getRs_dataRam_000();
        let x_9 = (victimLine_000);
        victims_000 <= update (x_6, x_7, Struct25 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct24 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_000 <= Struct24 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct29 x_10 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(3))'(3'h0))) begin
            let x_11 <- putRq_infoRam_000_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h1))) begin
            let x_13 <- putRq_infoRam_000_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h2))) begin
            let x_15 <- putRq_infoRam_000_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h3))) begin
            let x_17 <- putRq_infoRam_000_3(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h4))) begin
            let x_19 <- putRq_infoRam_000_4(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h5))) begin
            let x_21 <- putRq_infoRam_000_5(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h6))) begin
            let x_23 <- putRq_infoRam_000_6(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h7))) begin
            let x_25 <- putRq_infoRam_000_7(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_28 <- putRq_dataRam_000(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_000_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_000);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_000);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_000);
        Struct25 x_4 = ((x_3)[(Bit#(3))'(3'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_000 <= (Bit#(2))'(2'h3);
        readLine_000 <= (x_4).victim_line;

        end else begin

            Struct25 x_5 = ((x_3)[(Bit#(3))'(3'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_000 <= (Bit#(2))'(2'h3);
                readLine_000 <= (x_5).victim_line;

            end else begin

                Struct25 x_6 = ((x_3)[(Bit#(3))'(3'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_000 <= (Bit#(2))'(2'h3);
                    readLine_000 <= (x_6).victim_line;

                end else begin

                    Struct25 x_7 = ((x_3)[(Bit#(3))'(3'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_000 <= (Bit#(2))'(2'h3);
                        readLine_000 <= (x_7).victim_line;

                    end else begin

                        Struct25 x_8 = ((x_3)[(Bit#(3))'(3'h4)]);
                        if (((x_8).victim_valid) &&
                        ((((x_8).victim_line).addr) == (x_0))) begin

                            readStage_000 <= (Bit#(2))'(2'h3);
                            readLine_000 <= (x_8).victim_line;

                        end else begin

                            Struct25 x_9 = ((x_3)[(Bit#(3))'(3'h5)]);
                            if (((x_9).victim_valid) &&
                            ((((x_9).victim_line).addr) == (x_0))) begin

                                readStage_000 <= (Bit#(2))'(2'h3);

                                readLine_000 <= (x_9).victim_line;

                            end else begin

                                Struct25 x_10 = ((x_3)[(Bit#(3))'(3'h6)]);
                                if (((x_10).victim_valid) &&
                                ((((x_10).victim_line).addr) == (x_0))) begin

                                    readStage_000 <= (Bit#(2))'(2'h3);

                                    readLine_000 <= (x_10).victim_line;

                                end else begin

                                    Struct25 x_11 = ((x_3)[(Bit#(3))'(3'h7)]);

                                    if (((x_11).victim_valid) &&
                                    ((((x_11).victim_line).addr) == (x_0)))
                                    begin

                                        readStage_000 <= (Bit#(2))'(2'h3);

                                        readLine_000 <= (x_11).victim_line;

                                    end else begin

                                        readStage_000 <= (Bit#(2))'(2'h1);

                                        readAddr_000 <= x_0;
                                        Bit#(8) x_12 = ((x_0)[10:3]);
                                        Struct29 x_13 = (Struct29 {write :
                                        (Bool)'(False), addr : x_12, datain :
                                        (Struct26)'(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                                        let x_14 <-
                                        putRq_infoRam_000_0(x_13);
                                        let x_15 <-
                                        putRq_infoRam_000_1(x_13);
                                        let x_16 <-
                                        putRq_infoRam_000_2(x_13);
                                        let x_17 <-
                                        putRq_infoRam_000_3(x_13);
                                        let x_18 <-
                                        putRq_infoRam_000_4(x_13);
                                        let x_19 <-
                                        putRq_infoRam_000_5(x_13);
                                        let x_20 <-
                                        putRq_infoRam_000_6(x_13);
                                        let x_21 <-
                                        putRq_infoRam_000_7(x_13);

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_000_readRs ();
        let x_1 = (readStage_000);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_000 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_000);
        return x_2;
    endmethod

    method Action cache_000_writeRq (Struct24 x_0);
        let x_1 = (readStage_000);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_000);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_000);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct25 x_5 = ((x_3)[(Bit#(3))'(3'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct24 x_6 = (Struct24 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_000 <= x_6;
            victims_000 <= update (x_3, (Bit#(3))'(3'h0), Struct25
            {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h0), victim_line :
            x_6});

        end else begin

            Struct25 x_7 = ((x_3)[(Bit#(3))'(3'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct24 x_8 = (Struct24 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_000 <= x_8;
                victims_000 <= update (x_3, (Bit#(3))'(3'h1), Struct25
                {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h1),
                victim_line : x_8});

            end else begin

                Struct25 x_9 = ((x_3)[(Bit#(3))'(3'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct24 x_10 = (Struct24 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_000 <= x_10;
                    victims_000 <= update (x_3, (Bit#(3))'(3'h2), Struct25
                    {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h2),
                    victim_line : x_10});

                end else begin

                    Struct25 x_11 = ((x_3)[(Bit#(3))'(3'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct24 x_12 = (Struct24 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_000 <= x_12;
                        victims_000 <= update (x_3, (Bit#(3))'(3'h3),
                        Struct25 {victim_valid : x_4, victim_idx :
                        (Bit#(3))'(3'h3), victim_line : x_12});

                    end else begin

                        Struct25 x_13 = ((x_3)[(Bit#(3))'(3'h4)]);
                        if (((x_13).victim_valid) &&
                        ((((x_13).victim_line).addr) == ((x_0).addr))) begin

                            Struct24 x_14 = (Struct24 {addr : (x_0).addr,
                            info_hit : (Bool)'(False), info_way :
                            (x_0).info_way, info_write : (x_0).info_write,
                            info : (x_0).info, value_write :
                            (x_0).value_write, value : (x_0).value});

                            writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                            ((Bit#(3))'(3'h1)));
                            writeLine_000 <= x_14;
                            victims_000 <= update (x_3, (Bit#(3))'(3'h4),
                            Struct25 {victim_valid : x_4, victim_idx :
                            (Bit#(3))'(3'h4), victim_line : x_14});

                        end else begin

                            Struct25 x_15 = ((x_3)[(Bit#(3))'(3'h5)]);
                            if (((x_15).victim_valid) &&
                            ((((x_15).victim_line).addr) == ((x_0).addr)))
                            begin

                                Struct24 x_16 = (Struct24 {addr : (x_0).addr,
                                info_hit : (Bool)'(False), info_way :
                                (x_0).info_way, info_write :
                                (x_0).info_write, info : (x_0).info,
                                value_write : (x_0).value_write, value :
                                (x_0).value});
                                writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                                ((Bit#(3))'(3'h1)));
                                writeLine_000 <= x_16;
                                victims_000 <= update (x_3, (Bit#(3))'(3'h5),
                                Struct25 {victim_valid : x_4, victim_idx :
                                (Bit#(3))'(3'h5), victim_line : x_16});

                            end else begin

                                Struct25 x_17 = ((x_3)[(Bit#(3))'(3'h6)]);
                                if (((x_17).victim_valid) &&
                                ((((x_17).victim_line).addr) ==
                                ((x_0).addr))) begin

                                    Struct24 x_18 = (Struct24 {addr :
                                    (x_0).addr, info_hit : (Bool)'(False),
                                    info_way : (x_0).info_way, info_write :
                                    (x_0).info_write, info : (x_0).info,
                                    value_write : (x_0).value_write, value :
                                    (x_0).value});
                                    writeStage_000 <= (x_4 ?
                                    ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h1)));

                                    writeLine_000 <= x_18;
                                    victims_000 <= update (x_3,
                                    (Bit#(3))'(3'h6), Struct25 {victim_valid
                                    : x_4, victim_idx : (Bit#(3))'(3'h6),
                                    victim_line : x_18});

                                end else begin

                                    Struct25 x_19 = ((x_3)[(Bit#(3))'(3'h7)]);

                                    if (((x_19).victim_valid) &&
                                    ((((x_19).victim_line).addr) ==
                                    ((x_0).addr))) begin

                                        Struct24 x_20 = (Struct24 {addr :
                                        (x_0).addr, info_hit :
                                        (Bool)'(False), info_way :
                                        (x_0).info_way, info_write :
                                        (x_0).info_write, info : (x_0).info,
                                        value_write : (x_0).value_write,
                                        value : (x_0).value});
                                        writeStage_000 <= (x_4 ?
                                        ((Bit#(3))'(3'h7)) :
                                        ((Bit#(3))'(3'h1)));
                                        writeLine_000 <= x_20;
                                        victims_000 <= update (x_3,
                                        (Bit#(3))'(3'h7), Struct25
                                        {victim_valid : x_4, victim_idx :
                                        (Bit#(3))'(3'h7), victim_line :
                                        x_20});

                                    end else begin

                                        writeStage_000 <= (Bit#(3))'(3'h1);

                                        writeLine_000 <= x_0;

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_000_writeRs ();
        let x_1 = (writeStage_000);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_000 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_000);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_000_hasVictimSlot ();
        let x_1 = (victims_000);
        Bool x_2 = ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) ||
        (((x_1)[(Bit#(3))'(3'h0)]).victim_valid))))))));
        return x_2;
    endmethod

    method ActionValue#(Struct24) cache_000_getVictim ();
        let x_1 = (victims_000);
        when ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) ||
        (((x_1)[(Bit#(3))'(3'h0)]).victim_valid))))))), noAction);
        Struct24 x_2 = ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h7)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h6)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h5)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h4)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h3)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h2)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h1)]).victim_line) :
        (((x_1)[(Bit#(3))'(3'h0)]).victim_line)))))))))))))));
        return x_2;
    endmethod

    method Action cache_000_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_000);
        Struct25 x_2 = ((x_1)[(Bit#(3))'(3'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_000 <= update (x_1, (Bit#(3))'(3'h0),
            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct25 x_3 = ((x_1)[(Bit#(3))'(3'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_000 <= update (x_1, (Bit#(3))'(3'h1),
                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct25 x_4 = ((x_1)[(Bit#(3))'(3'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_000 <= update (x_1, (Bit#(3))'(3'h2),
                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct25 x_5 = ((x_1)[(Bit#(3))'(3'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_000 <= update (x_1, (Bit#(3))'(3'h3),
                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                        Struct25 x_6 = ((x_1)[(Bit#(3))'(3'h4)]);
                        if (((x_6).victim_valid) &&
                        ((((x_6).victim_line).addr) == (x_0))) begin

                            victims_000 <= update (x_1, (Bit#(3))'(3'h4),
                            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                        end else begin

                            Struct25 x_7 = ((x_1)[(Bit#(3))'(3'h5)]);
                            if (((x_7).victim_valid) &&
                            ((((x_7).victim_line).addr) == (x_0))) begin

                                victims_000 <= update (x_1, (Bit#(3))'(3'h5),
                                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                            end else begin

                                Struct25 x_8 = ((x_1)[(Bit#(3))'(3'h6)]);
                                if (((x_8).victim_valid) &&
                                ((((x_8).victim_line).addr) == (x_0))) begin

                                    victims_000 <= update (x_1,
                                    (Bit#(3))'(3'h6),
                                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                                end else begin

                                    Struct25 x_9 = ((x_1)[(Bit#(3))'(3'h7)]);

                                    if (((x_9).victim_valid) &&
                                    ((((x_9).victim_line).addr) == (x_0)))
                                    begin

                                        victims_000 <= update (x_1,
                                        (Bit#(3))'(3'h7),
                                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                                    end else begin

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

endmodule

interface Module136;
    method Action makeEnq_parentChildren000 (Struct10 x_0);
    method Action broadcast_parentChildren000 (Struct13 x_0);

endinterface


module mkModule136#(function Action enq_fifo00002(Struct2 _),
  function Action enq_fifo00012(Struct2 _),
  function Action enq_fifo00022(Struct2 _),
  function Action enq_fifo00032(Struct2 _),
  function Action enq_fifo0001(Struct2 _),
  function Action enq_fifo0000(Struct2 _)) (Module136);

    // No rules in this module

    method Action makeEnq_parentChildren000 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo0000((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo0001((x_0).enq_msg);

            end else begin

                Bit#(2) x_3 = ((x_0).enq_ch_idx);
                Struct2 x_4 = ((x_0).enq_msg);
                if ((x_3) == ((Bit#(2))'(2'h3))) begin
                let x_5 <- enq_fifo00032(x_4);

                end else begin

                    if ((x_3) == ((Bit#(2))'(2'h2))) begin
                    let x_6 <- enq_fifo00022(x_4);

                    end else begin

                        if ((x_3) == ((Bit#(2))'(2'h1))) begin
                        let x_7 <- enq_fifo00012(x_4);

                        end else begin

                            if ((x_3) == ((Bit#(2))'(2'h0))) begin
                            let x_8 <- enq_fifo00002(x_4);

                            end else begin

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method Action broadcast_parentChildren000 (Struct13 x_0);
        Bit#(4) x_1 = ((x_0).cs_inds);
        Struct2 x_2 = ((x_0).cs_msg);
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == (x_1))
        begin
        let x_3 <- enq_fifo00032(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == (x_1))
        begin
        let x_5 <- enq_fifo00022(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == (x_1))
        begin
        let x_7 <- enq_fifo00012(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == (x_1))
        begin
        let x_9 <- enq_fifo00002(x_2);

        end else begin

        end

    endmethod

endmodule

interface Module137;
    method Action cache_0000_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0000_readRs ();
    method Action cache_0000_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0000_writeRs ();
    method ActionValue#(Bool) cache_0000_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0000_getVictim ();
    method Action cache_0000_removeVictim (Bit#(64) x_0);

endinterface


module mkModule137#(function Action putRq_infoRam_0000_3(Struct36 _),
  function Action putRq_infoRam_0000_2(Struct36 _),
  function Action putRq_infoRam_0000_1(Struct36 _),
  function Action putRq_infoRam_0000_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0000(),
  function Action putRq_dataRam_0000(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0000_3(),
  function ActionValue#(Struct33) getRs_infoRam_0000_2(),
  function ActionValue#(Struct33) getRs_infoRam_0000_1(),
  function ActionValue#(Struct33) getRs_infoRam_0000_0()) (Module137);
    Reg#(Bit#(2)) readStage_0000 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0000 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0000 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0000 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0000 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0000 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0000 <- mkReg(unpack(0));

    rule read_tagmatch_0000;
        let x_0 = (readStage_0000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0000);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0000_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0000_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0000_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0000_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0000 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0000 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0000(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0000 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0000;
        let x_0 = (readStage_0000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0000 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0000();
        let x_2 = (readLine_0000);
        readLine_0000 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0000;
        let x_0 = (writeStage_0000);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0000);
        when ((x_1).info_hit, noAction);
        writeStage_0000 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0000_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0000_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0000_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0000_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0000(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0000;
        let x_0 = (writeStage_0000);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0000);
        when (! ((x_1).info_hit), noAction);
        writeStage_0000 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0000_0(x_4);
        let x_6 <- putRq_infoRam_0000_1(x_4);
        let x_7 <- putRq_infoRam_0000_2(x_4);
        let x_8 <- putRq_infoRam_0000_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0000;
        let x_0 = (writeStage_0000);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0000 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0000_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0000_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0000_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0000_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0000);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0000 <= x_10;
        victimLine_0000 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0000(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0000;
        let x_0 = (writeStage_0000);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0000);
        writeStage_0000 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0000);
        let x_6 = (victims_0000);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0000();
        let x_9 = (victimLine_0000);
        victims_0000 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0000 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0000_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0000_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0000_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0000_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0000(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0000_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0000);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0000);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0000);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0000 <= (Bit#(2))'(2'h3);
            readLine_0000 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0000 <= (Bit#(2))'(2'h3);
                readLine_0000 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0000 <= (Bit#(2))'(2'h3);
                    readLine_0000 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0000 <= (Bit#(2))'(2'h3);
                        readLine_0000 <= (x_7).victim_line;

                    end else begin

                        readStage_0000 <= (Bit#(2))'(2'h1);
                        readAddr_0000 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0000_0(x_9);
                        let x_11 <- putRq_infoRam_0000_1(x_9);
                        let x_12 <- putRq_infoRam_0000_2(x_9);
                        let x_13 <- putRq_infoRam_0000_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0000_readRs ();
        let x_1 = (readStage_0000);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0000 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0000);
        return x_2;
    endmethod

    method Action cache_0000_writeRq (Struct31 x_0);
        let x_1 = (readStage_0000);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0000);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0000);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0000 <= x_6;
            victims_0000 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0000 <= x_8;
                victims_0000 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0000 <= x_10;
                    victims_0000 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0000 <= x_12;
                        victims_0000 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0000 <= (Bit#(3))'(3'h1);
                        writeLine_0000 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0000_writeRs ();
        let x_1 = (writeStage_0000);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0000 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0000);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0000_hasVictimSlot ();
        let x_1 = (victims_0000);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0000_getVictim ();
        let x_1 = (victims_0000);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0000_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0000);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0000 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0000 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0000 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0000 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module138; method Action makeEnq_parentChildren0000 (Struct10 x_0);

endinterface


module mkModule138#(function Action enq_fifo000002(Struct2 _),
  function Action enq_fifo00001(Struct2 _),
  function Action enq_fifo00000(Struct2 _)) (Module138);

    // No rules in this module

    method Action makeEnq_parentChildren0000 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00000((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00001((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo000002(x_3);

            end

        end

    endmethod

endmodule

interface Module139;
    method Action cache_0001_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0001_readRs ();
    method Action cache_0001_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0001_writeRs ();
    method ActionValue#(Bool) cache_0001_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0001_getVictim ();
    method Action cache_0001_removeVictim (Bit#(64) x_0);

endinterface


module mkModule139#(function Action putRq_infoRam_0001_3(Struct36 _),
  function Action putRq_infoRam_0001_2(Struct36 _),
  function Action putRq_infoRam_0001_1(Struct36 _),
  function Action putRq_infoRam_0001_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0001(),
  function Action putRq_dataRam_0001(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0001_3(),
  function ActionValue#(Struct33) getRs_infoRam_0001_2(),
  function ActionValue#(Struct33) getRs_infoRam_0001_1(),
  function ActionValue#(Struct33) getRs_infoRam_0001_0()) (Module139);
    Reg#(Bit#(2)) readStage_0001 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0001 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0001 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0001 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0001 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0001 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0001 <- mkReg(unpack(0));

    rule read_tagmatch_0001;
        let x_0 = (readStage_0001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0001);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0001_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0001_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0001_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0001_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0001 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0001 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0001(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0001 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0001;
        let x_0 = (readStage_0001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0001 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0001();
        let x_2 = (readLine_0001);
        readLine_0001 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0001;
        let x_0 = (writeStage_0001);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0001);
        when ((x_1).info_hit, noAction);
        writeStage_0001 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0001_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0001_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0001_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0001_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0001(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0001;
        let x_0 = (writeStage_0001);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0001);
        when (! ((x_1).info_hit), noAction);
        writeStage_0001 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0001_0(x_4);
        let x_6 <- putRq_infoRam_0001_1(x_4);
        let x_7 <- putRq_infoRam_0001_2(x_4);
        let x_8 <- putRq_infoRam_0001_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0001;
        let x_0 = (writeStage_0001);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0001 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0001_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0001_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0001_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0001_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0001);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0001 <= x_10;
        victimLine_0001 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0001(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0001;
        let x_0 = (writeStage_0001);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0001);
        writeStage_0001 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0001);
        let x_6 = (victims_0001);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0001();
        let x_9 = (victimLine_0001);
        victims_0001 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0001 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0001_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0001_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0001_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0001_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0001(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0001_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0001);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0001);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0001);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0001 <= (Bit#(2))'(2'h3);
            readLine_0001 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0001 <= (Bit#(2))'(2'h3);
                readLine_0001 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0001 <= (Bit#(2))'(2'h3);
                    readLine_0001 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0001 <= (Bit#(2))'(2'h3);
                        readLine_0001 <= (x_7).victim_line;

                    end else begin

                        readStage_0001 <= (Bit#(2))'(2'h1);
                        readAddr_0001 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0001_0(x_9);
                        let x_11 <- putRq_infoRam_0001_1(x_9);
                        let x_12 <- putRq_infoRam_0001_2(x_9);
                        let x_13 <- putRq_infoRam_0001_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0001_readRs ();
        let x_1 = (readStage_0001);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0001 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0001);
        return x_2;
    endmethod

    method Action cache_0001_writeRq (Struct31 x_0);
        let x_1 = (readStage_0001);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0001);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0001);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0001 <= x_6;
            victims_0001 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0001 <= x_8;
                victims_0001 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0001 <= x_10;
                    victims_0001 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0001 <= x_12;
                        victims_0001 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0001 <= (Bit#(3))'(3'h1);
                        writeLine_0001 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0001_writeRs ();
        let x_1 = (writeStage_0001);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0001 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0001);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0001_hasVictimSlot ();
        let x_1 = (victims_0001);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0001_getVictim ();
        let x_1 = (victims_0001);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0001_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0001);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0001 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0001 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0001 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0001 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module140; method Action makeEnq_parentChildren0001 (Struct10 x_0);

endinterface


module mkModule140#(function Action enq_fifo000102(Struct2 _),
  function Action enq_fifo00011(Struct2 _),
  function Action enq_fifo00010(Struct2 _)) (Module140);

    // No rules in this module

    method Action makeEnq_parentChildren0001 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00010((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00011((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo000102(x_3);

            end

        end

    endmethod

endmodule

interface Module141;
    method Action cache_0002_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0002_readRs ();
    method Action cache_0002_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0002_writeRs ();
    method ActionValue#(Bool) cache_0002_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0002_getVictim ();
    method Action cache_0002_removeVictim (Bit#(64) x_0);

endinterface


module mkModule141#(function Action putRq_infoRam_0002_3(Struct36 _),
  function Action putRq_infoRam_0002_2(Struct36 _),
  function Action putRq_infoRam_0002_1(Struct36 _),
  function Action putRq_infoRam_0002_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0002(),
  function Action putRq_dataRam_0002(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0002_3(),
  function ActionValue#(Struct33) getRs_infoRam_0002_2(),
  function ActionValue#(Struct33) getRs_infoRam_0002_1(),
  function ActionValue#(Struct33) getRs_infoRam_0002_0()) (Module141);
    Reg#(Bit#(2)) readStage_0002 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0002 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0002 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0002 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0002 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0002 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0002 <- mkReg(unpack(0));

    rule read_tagmatch_0002;
        let x_0 = (readStage_0002);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0002);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0002_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0002_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0002_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0002_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0002 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0002 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0002(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0002 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0002;
        let x_0 = (readStage_0002);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0002 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0002();
        let x_2 = (readLine_0002);
        readLine_0002 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0002;
        let x_0 = (writeStage_0002);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0002);
        when ((x_1).info_hit, noAction);
        writeStage_0002 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0002_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0002_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0002_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0002_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0002(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0002;
        let x_0 = (writeStage_0002);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0002);
        when (! ((x_1).info_hit), noAction);
        writeStage_0002 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0002_0(x_4);
        let x_6 <- putRq_infoRam_0002_1(x_4);
        let x_7 <- putRq_infoRam_0002_2(x_4);
        let x_8 <- putRq_infoRam_0002_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0002;
        let x_0 = (writeStage_0002);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0002 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0002_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0002_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0002_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0002_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0002);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0002 <= x_10;
        victimLine_0002 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0002(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0002;
        let x_0 = (writeStage_0002);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0002);
        writeStage_0002 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0002);
        let x_6 = (victims_0002);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0002();
        let x_9 = (victimLine_0002);
        victims_0002 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0002 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0002_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0002_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0002_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0002_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0002(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0002_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0002);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0002);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0002);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0002 <= (Bit#(2))'(2'h3);
            readLine_0002 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0002 <= (Bit#(2))'(2'h3);
                readLine_0002 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0002 <= (Bit#(2))'(2'h3);
                    readLine_0002 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0002 <= (Bit#(2))'(2'h3);
                        readLine_0002 <= (x_7).victim_line;

                    end else begin

                        readStage_0002 <= (Bit#(2))'(2'h1);
                        readAddr_0002 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0002_0(x_9);
                        let x_11 <- putRq_infoRam_0002_1(x_9);
                        let x_12 <- putRq_infoRam_0002_2(x_9);
                        let x_13 <- putRq_infoRam_0002_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0002_readRs ();
        let x_1 = (readStage_0002);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0002 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0002);
        return x_2;
    endmethod

    method Action cache_0002_writeRq (Struct31 x_0);
        let x_1 = (readStage_0002);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0002);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0002);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0002 <= x_6;
            victims_0002 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0002 <= x_8;
                victims_0002 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0002 <= x_10;
                    victims_0002 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0002 <= x_12;
                        victims_0002 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0002 <= (Bit#(3))'(3'h1);
                        writeLine_0002 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0002_writeRs ();
        let x_1 = (writeStage_0002);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0002 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0002);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0002_hasVictimSlot ();
        let x_1 = (victims_0002);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0002_getVictim ();
        let x_1 = (victims_0002);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0002_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0002);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0002 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0002 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0002 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0002 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module142; method Action makeEnq_parentChildren0002 (Struct10 x_0);

endinterface


module mkModule142#(function Action enq_fifo000202(Struct2 _),
  function Action enq_fifo00021(Struct2 _),
  function Action enq_fifo00020(Struct2 _)) (Module142);

    // No rules in this module

    method Action makeEnq_parentChildren0002 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00020((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00021((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo000202(x_3);

            end

        end

    endmethod

endmodule

interface Module143;
    method Action cache_0003_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0003_readRs ();
    method Action cache_0003_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0003_writeRs ();
    method ActionValue#(Bool) cache_0003_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0003_getVictim ();
    method Action cache_0003_removeVictim (Bit#(64) x_0);

endinterface


module mkModule143#(function Action putRq_infoRam_0003_3(Struct36 _),
  function Action putRq_infoRam_0003_2(Struct36 _),
  function Action putRq_infoRam_0003_1(Struct36 _),
  function Action putRq_infoRam_0003_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0003(),
  function Action putRq_dataRam_0003(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0003_3(),
  function ActionValue#(Struct33) getRs_infoRam_0003_2(),
  function ActionValue#(Struct33) getRs_infoRam_0003_1(),
  function ActionValue#(Struct33) getRs_infoRam_0003_0()) (Module143);
    Reg#(Bit#(2)) readStage_0003 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0003 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0003 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0003 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0003 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0003 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0003 <- mkReg(unpack(0));

    rule read_tagmatch_0003;
        let x_0 = (readStage_0003);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0003);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0003_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0003_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0003_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0003_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0003 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0003 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0003(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0003 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0003;
        let x_0 = (readStage_0003);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0003 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0003();
        let x_2 = (readLine_0003);
        readLine_0003 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0003;
        let x_0 = (writeStage_0003);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0003);
        when ((x_1).info_hit, noAction);
        writeStage_0003 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0003_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0003_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0003_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0003_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0003(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0003;
        let x_0 = (writeStage_0003);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0003);
        when (! ((x_1).info_hit), noAction);
        writeStage_0003 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0003_0(x_4);
        let x_6 <- putRq_infoRam_0003_1(x_4);
        let x_7 <- putRq_infoRam_0003_2(x_4);
        let x_8 <- putRq_infoRam_0003_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0003;
        let x_0 = (writeStage_0003);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0003 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0003_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0003_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0003_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0003_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0003);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0003 <= x_10;
        victimLine_0003 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0003(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0003;
        let x_0 = (writeStage_0003);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0003);
        writeStage_0003 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0003);
        let x_6 = (victims_0003);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0003();
        let x_9 = (victimLine_0003);
        victims_0003 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0003 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0003_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0003_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0003_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0003_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0003(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0003_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0003);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0003);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0003);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0003 <= (Bit#(2))'(2'h3);
            readLine_0003 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0003 <= (Bit#(2))'(2'h3);
                readLine_0003 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0003 <= (Bit#(2))'(2'h3);
                    readLine_0003 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0003 <= (Bit#(2))'(2'h3);
                        readLine_0003 <= (x_7).victim_line;

                    end else begin

                        readStage_0003 <= (Bit#(2))'(2'h1);
                        readAddr_0003 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0003_0(x_9);
                        let x_11 <- putRq_infoRam_0003_1(x_9);
                        let x_12 <- putRq_infoRam_0003_2(x_9);
                        let x_13 <- putRq_infoRam_0003_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0003_readRs ();
        let x_1 = (readStage_0003);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0003 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0003);
        return x_2;
    endmethod

    method Action cache_0003_writeRq (Struct31 x_0);
        let x_1 = (readStage_0003);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0003);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0003);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0003 <= x_6;
            victims_0003 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0003 <= x_8;
                victims_0003 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0003 <= x_10;
                    victims_0003 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0003 <= x_12;
                        victims_0003 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0003 <= (Bit#(3))'(3'h1);
                        writeLine_0003 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0003_writeRs ();
        let x_1 = (writeStage_0003);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0003 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0003);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0003_hasVictimSlot ();
        let x_1 = (victims_0003);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0003_getVictim ();
        let x_1 = (victims_0003);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0003_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0003);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0003 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0003 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0003 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0003 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module144; method Action makeEnq_parentChildren0003 (Struct10 x_0);

endinterface


module mkModule144#(function Action enq_fifo000302(Struct2 _),
  function Action enq_fifo00031(Struct2 _),
  function Action enq_fifo00030(Struct2 _)) (Module144);

    // No rules in this module

    method Action makeEnq_parentChildren0003 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00030((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00031((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo000302(x_3);

            end

        end

    endmethod

endmodule

interface Module145;
    method Action cache_001_readRq (Bit#(64) x_0);
    method ActionValue#(Struct24) cache_001_readRs ();
    method Action cache_001_writeRq (Struct24 x_0);
    method ActionValue#(Struct24) cache_001_writeRs ();
    method ActionValue#(Bool) cache_001_hasVictimSlot ();
    method ActionValue#(Struct24) cache_001_getVictim ();
    method Action cache_001_removeVictim (Bit#(64) x_0);

endinterface


module mkModule145#(function Action putRq_infoRam_001_7(Struct29 _),
  function Action putRq_infoRam_001_6(Struct29 _),
  function Action putRq_infoRam_001_5(Struct29 _),
  function Action putRq_infoRam_001_4(Struct29 _),
  function Action putRq_infoRam_001_3(Struct29 _),
  function Action putRq_infoRam_001_2(Struct29 _),
  function Action putRq_infoRam_001_1(Struct29 _),
  function Action putRq_infoRam_001_0(Struct29 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_001(),
  function Action putRq_dataRam_001(Struct28 _),
  function ActionValue#(Struct26) getRs_infoRam_001_7(),
  function ActionValue#(Struct26) getRs_infoRam_001_6(),
  function ActionValue#(Struct26) getRs_infoRam_001_5(),
  function ActionValue#(Struct26) getRs_infoRam_001_4(),
  function ActionValue#(Struct26) getRs_infoRam_001_3(),
  function ActionValue#(Struct26) getRs_infoRam_001_2(),
  function ActionValue#(Struct26) getRs_infoRam_001_1(),
  function ActionValue#(Struct26) getRs_infoRam_001_0()) (Module145);
    Reg#(Bit#(2)) readStage_001 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_001 <- mkReg(unpack(0));
    Reg#(Struct24) readLine_001 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_001 <- mkReg(unpack(0));
    Reg#(Struct24) writeLine_001 <- mkReg(unpack(0));
    Reg#(Vector#(8, Struct25)) victims_001 <- mkReg(unpack(0));
    Reg#(Struct24) victimLine_001 <- mkReg(unpack(0));
    Reg#(Bit#(3)) victimWay_001 <- mkReg(unpack(0));

    rule read_tagmatch_001;
        let x_0 = (readStage_001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_001);
        Bit#(53) x_2 = ((x_1)[63:11]);
        Bit#(8) x_3 = ((x_1)[10:3]);
        Vector#(8, Struct26) x_4 =
        ((Vector#(8, Struct26))'(vec(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_001_0();
        Vector#(8, Struct26) x_6 = (update (x_4, (Bit#(3))'(3'h0), x_5));
        let x_7 <- getRs_infoRam_001_1();
        Vector#(8, Struct26) x_8 = (update (x_6, (Bit#(3))'(3'h1), x_7));
        let x_9 <- getRs_infoRam_001_2();
        Vector#(8, Struct26) x_10 = (update (x_8, (Bit#(3))'(3'h2), x_9));
        let x_11 <- getRs_infoRam_001_3();
        Vector#(8, Struct26) x_12 = (update (x_10, (Bit#(3))'(3'h3), x_11));

        let x_13 <- getRs_infoRam_001_4();
        Vector#(8, Struct26) x_14 = (update (x_12, (Bit#(3))'(3'h4), x_13));

        let x_15 <- getRs_infoRam_001_5();
        Vector#(8, Struct26) x_16 = (update (x_14, (Bit#(3))'(3'h5), x_15));

        let x_17 <- getRs_infoRam_001_6();
        Vector#(8, Struct26) x_18 = (update (x_16, (Bit#(3))'(3'h6), x_17));

        let x_19 <- getRs_infoRam_001_7();
        Vector#(8, Struct26) x_20 = (update (x_18, (Bit#(3))'(3'h7), x_19));

        Struct27 x_21 = (((((x_20)[(Bit#(3))'(3'h0)]).tag) == (x_2) ?
        (Struct27 {tm_hit : (Bool)'(True), tm_way : (Bit#(3))'(3'h0),
        tm_value : ((x_20)[(Bit#(3))'(3'h0)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h1)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h1), tm_value :
        ((x_20)[(Bit#(3))'(3'h1)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h2)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h2), tm_value :
        ((x_20)[(Bit#(3))'(3'h2)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h3)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h3), tm_value :
        ((x_20)[(Bit#(3))'(3'h3)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h4)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h4), tm_value :
        ((x_20)[(Bit#(3))'(3'h4)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h5)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h5), tm_value :
        ((x_20)[(Bit#(3))'(3'h5)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h6)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h6), tm_value :
        ((x_20)[(Bit#(3))'(3'h6)]).value}) :
        (((((x_20)[(Bit#(3))'(3'h7)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(3))'(3'h7), tm_value :
        ((x_20)[(Bit#(3))'(3'h7)]).value}) :
        ((Struct27)'(Struct27 {tm_hit: False, tm_way: 3'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))))))))))));

        readLine_001 <= Struct24 {addr : x_1, info_hit : (x_21).tm_hit,
        info_way : (x_21).tm_way, info_write : (Bool)'(False), info :
        (x_21).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_21).tm_hit) begin

            readStage_001 <= (Bit#(2))'(2'h2);
            let x_22 <- putRq_dataRam_001(Struct28 {write : (Bool)'(False),
            addr : {(x_3),((x_21).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_001 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_001;
        let x_0 = (readStage_001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_001 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_001();
        let x_2 = (readLine_001);
        readLine_001 <= Struct24 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_001);
        when ((x_1).info_hit, noAction);
        writeStage_001 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(53) x_3 = ((x_2)[63:11]);
        Bit#(8) x_4 = ((x_2)[10:3]);
        Bit#(3) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct29 x_6 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(3))'(3'h0))) begin
            let x_7 <- putRq_infoRam_001_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h1))) begin
            let x_9 <- putRq_infoRam_001_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h2))) begin
            let x_11 <- putRq_infoRam_001_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h3))) begin
            let x_13 <- putRq_infoRam_001_3(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h4))) begin
            let x_15 <- putRq_infoRam_001_4(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h5))) begin
            let x_17 <- putRq_infoRam_001_5(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h6))) begin
            let x_19 <- putRq_infoRam_001_6(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h7))) begin
            let x_21 <- putRq_infoRam_001_7(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_24 <- putRq_dataRam_001(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_001);
        when (! ((x_1).info_hit), noAction);
        writeStage_001 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(8) x_3 = ((x_2)[10:3]);
        Struct29 x_4 = (Struct29 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct26)'(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_001_0(x_4);
        let x_6 <- putRq_infoRam_001_1(x_4);
        let x_7 <- putRq_infoRam_001_2(x_4);
        let x_8 <- putRq_infoRam_001_3(x_4);
        let x_9 <- putRq_infoRam_001_4(x_4);
        let x_10 <- putRq_infoRam_001_5(x_4);
        let x_11 <- putRq_infoRam_001_6(x_4);
        let x_12 <- putRq_infoRam_001_7(x_4);

    endrule

    rule write_info_miss_rep_rs_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_001 <= (Bit#(3))'(3'h3);
        Vector#(8, Struct26) x_1 =
        ((Vector#(8, Struct26))'(vec(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_001_0();
        Vector#(8, Struct26) x_3 = (update (x_1, (Bit#(3))'(3'h0), x_2));
        let x_4 <- getRs_infoRam_001_1();
        Vector#(8, Struct26) x_5 = (update (x_3, (Bit#(3))'(3'h1), x_4));
        let x_6 <- getRs_infoRam_001_2();
        Vector#(8, Struct26) x_7 = (update (x_5, (Bit#(3))'(3'h2), x_6));
        let x_8 <- getRs_infoRam_001_3();
        Vector#(8, Struct26) x_9 = (update (x_7, (Bit#(3))'(3'h3), x_8));
        let x_10 <- getRs_infoRam_001_4();
        Vector#(8, Struct26) x_11 = (update (x_9, (Bit#(3))'(3'h4), x_10));

        let x_12 <- getRs_infoRam_001_5();
        Vector#(8, Struct26) x_13 = (update (x_11, (Bit#(3))'(3'h5), x_12));

        let x_14 <- getRs_infoRam_001_6();
        Vector#(8, Struct26) x_15 = (update (x_13, (Bit#(3))'(3'h6), x_14));

        let x_16 <- getRs_infoRam_001_7();
        Vector#(8, Struct26) x_17 = (update (x_15, (Bit#(3))'(3'h7), x_16));

        Bit#(3) x_18 = ((((((x_17)[(Bit#(3))'(3'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h0)) :
        ((((((x_17)[(Bit#(3))'(3'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h1)) :
        ((((((x_17)[(Bit#(3))'(3'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h2)) :
        ((((((x_17)[(Bit#(3))'(3'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h3)) :
        ((((((x_17)[(Bit#(3))'(3'h4)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h4)) :
        ((((((x_17)[(Bit#(3))'(3'h5)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h5)) :
        ((((((x_17)[(Bit#(3))'(3'h6)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h6)) :
        ((((((x_17)[(Bit#(3))'(3'h7)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(3))'(3'h7)) :
        ((Bit#(3))'(3'h0))))))))))))))))));
        let x_19 = (writeLine_001);
        Bit#(64) x_20 = ((x_19).addr);
        Bit#(8) x_21 = ((x_20)[10:3]);
        Struct26 x_22 = ((x_17)[x_18]);
        Bit#(53) x_23 = ((x_22).tag);
        Struct4 x_24 = ((x_22).value);
        victimWay_001 <= x_18;
        victimLine_001 <= Struct24 {addr :
        {(x_23),({(x_21),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(3))'(3'h0), info_write : (Bool)'(False), info :
        x_24, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_25 <- putRq_dataRam_001(Struct28 {write : (Bool)'(False), addr
        : {(x_21),(x_18)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_001);
        writeStage_001 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(53) x_3 = ((x_2)[63:11]);
        Bit#(8) x_4 = ((x_2)[10:3]);
        let x_5 = (victimWay_001);
        let x_6 = (victims_001);
        when ((! (((x_6)[(Bit#(3))'(3'h7)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h6)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h5)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h4)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(3))'(3'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(3))'(3'h0)]).victim_valid)))))))), noAction);
        Bit#(3) x_7 = ((((x_6)[(Bit#(3))'(3'h7)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h6)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h5)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h4)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h3)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h2)]).victim_valid ?
        ((((x_6)[(Bit#(3))'(3'h1)]).victim_valid ? ((Bit#(3))'(3'h0)) :
        ((Bit#(3))'(3'h1)))) : ((Bit#(3))'(3'h2)))) : ((Bit#(3))'(3'h3)))) :
        ((Bit#(3))'(3'h4)))) : ((Bit#(3))'(3'h5)))) : ((Bit#(3))'(3'h6)))) :
        ((Bit#(3))'(3'h7))));
        let x_8 <- getRs_dataRam_001();
        let x_9 = (victimLine_001);
        victims_001 <= update (x_6, x_7, Struct25 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct24 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_001 <= Struct24 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct29 x_10 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(3))'(3'h0))) begin
            let x_11 <- putRq_infoRam_001_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h1))) begin
            let x_13 <- putRq_infoRam_001_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h2))) begin
            let x_15 <- putRq_infoRam_001_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h3))) begin
            let x_17 <- putRq_infoRam_001_3(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h4))) begin
            let x_19 <- putRq_infoRam_001_4(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h5))) begin
            let x_21 <- putRq_infoRam_001_5(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h6))) begin
            let x_23 <- putRq_infoRam_001_6(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(3))'(3'h7))) begin
            let x_25 <- putRq_infoRam_001_7(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_28 <- putRq_dataRam_001(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_001_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_001);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_001);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_001);
        Struct25 x_4 = ((x_3)[(Bit#(3))'(3'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_001 <= (Bit#(2))'(2'h3);
        readLine_001 <= (x_4).victim_line;

        end else begin

            Struct25 x_5 = ((x_3)[(Bit#(3))'(3'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_001 <= (Bit#(2))'(2'h3);
                readLine_001 <= (x_5).victim_line;

            end else begin

                Struct25 x_6 = ((x_3)[(Bit#(3))'(3'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_001 <= (Bit#(2))'(2'h3);
                    readLine_001 <= (x_6).victim_line;

                end else begin

                    Struct25 x_7 = ((x_3)[(Bit#(3))'(3'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_001 <= (Bit#(2))'(2'h3);
                        readLine_001 <= (x_7).victim_line;

                    end else begin

                        Struct25 x_8 = ((x_3)[(Bit#(3))'(3'h4)]);
                        if (((x_8).victim_valid) &&
                        ((((x_8).victim_line).addr) == (x_0))) begin

                            readStage_001 <= (Bit#(2))'(2'h3);
                            readLine_001 <= (x_8).victim_line;

                        end else begin

                            Struct25 x_9 = ((x_3)[(Bit#(3))'(3'h5)]);
                            if (((x_9).victim_valid) &&
                            ((((x_9).victim_line).addr) == (x_0))) begin

                                readStage_001 <= (Bit#(2))'(2'h3);

                                readLine_001 <= (x_9).victim_line;

                            end else begin

                                Struct25 x_10 = ((x_3)[(Bit#(3))'(3'h6)]);
                                if (((x_10).victim_valid) &&
                                ((((x_10).victim_line).addr) == (x_0))) begin

                                    readStage_001 <= (Bit#(2))'(2'h3);

                                    readLine_001 <= (x_10).victim_line;

                                end else begin

                                    Struct25 x_11 = ((x_3)[(Bit#(3))'(3'h7)]);

                                    if (((x_11).victim_valid) &&
                                    ((((x_11).victim_line).addr) == (x_0)))
                                    begin

                                        readStage_001 <= (Bit#(2))'(2'h3);

                                        readLine_001 <= (x_11).victim_line;

                                    end else begin

                                        readStage_001 <= (Bit#(2))'(2'h1);

                                        readAddr_001 <= x_0;
                                        Bit#(8) x_12 = ((x_0)[10:3]);
                                        Struct29 x_13 = (Struct29 {write :
                                        (Bool)'(False), addr : x_12, datain :
                                        (Struct26)'(Struct26 {tag: 53'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                                        let x_14 <-
                                        putRq_infoRam_001_0(x_13);
                                        let x_15 <-
                                        putRq_infoRam_001_1(x_13);
                                        let x_16 <-
                                        putRq_infoRam_001_2(x_13);
                                        let x_17 <-
                                        putRq_infoRam_001_3(x_13);
                                        let x_18 <-
                                        putRq_infoRam_001_4(x_13);
                                        let x_19 <-
                                        putRq_infoRam_001_5(x_13);
                                        let x_20 <-
                                        putRq_infoRam_001_6(x_13);
                                        let x_21 <-
                                        putRq_infoRam_001_7(x_13);

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_001_readRs ();
        let x_1 = (readStage_001);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_001 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_001);
        return x_2;
    endmethod

    method Action cache_001_writeRq (Struct24 x_0);
        let x_1 = (readStage_001);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_001);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_001);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct25 x_5 = ((x_3)[(Bit#(3))'(3'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct24 x_6 = (Struct24 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_001 <= x_6;
            victims_001 <= update (x_3, (Bit#(3))'(3'h0), Struct25
            {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h0), victim_line :
            x_6});

        end else begin

            Struct25 x_7 = ((x_3)[(Bit#(3))'(3'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct24 x_8 = (Struct24 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_001 <= x_8;
                victims_001 <= update (x_3, (Bit#(3))'(3'h1), Struct25
                {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h1),
                victim_line : x_8});

            end else begin

                Struct25 x_9 = ((x_3)[(Bit#(3))'(3'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct24 x_10 = (Struct24 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_001 <= x_10;
                    victims_001 <= update (x_3, (Bit#(3))'(3'h2), Struct25
                    {victim_valid : x_4, victim_idx : (Bit#(3))'(3'h2),
                    victim_line : x_10});

                end else begin

                    Struct25 x_11 = ((x_3)[(Bit#(3))'(3'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct24 x_12 = (Struct24 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_001 <= x_12;
                        victims_001 <= update (x_3, (Bit#(3))'(3'h3),
                        Struct25 {victim_valid : x_4, victim_idx :
                        (Bit#(3))'(3'h3), victim_line : x_12});

                    end else begin

                        Struct25 x_13 = ((x_3)[(Bit#(3))'(3'h4)]);
                        if (((x_13).victim_valid) &&
                        ((((x_13).victim_line).addr) == ((x_0).addr))) begin

                            Struct24 x_14 = (Struct24 {addr : (x_0).addr,
                            info_hit : (Bool)'(False), info_way :
                            (x_0).info_way, info_write : (x_0).info_write,
                            info : (x_0).info, value_write :
                            (x_0).value_write, value : (x_0).value});

                            writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                            ((Bit#(3))'(3'h1)));
                            writeLine_001 <= x_14;
                            victims_001 <= update (x_3, (Bit#(3))'(3'h4),
                            Struct25 {victim_valid : x_4, victim_idx :
                            (Bit#(3))'(3'h4), victim_line : x_14});

                        end else begin

                            Struct25 x_15 = ((x_3)[(Bit#(3))'(3'h5)]);
                            if (((x_15).victim_valid) &&
                            ((((x_15).victim_line).addr) == ((x_0).addr)))
                            begin

                                Struct24 x_16 = (Struct24 {addr : (x_0).addr,
                                info_hit : (Bool)'(False), info_way :
                                (x_0).info_way, info_write :
                                (x_0).info_write, info : (x_0).info,
                                value_write : (x_0).value_write, value :
                                (x_0).value});
                                writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                                ((Bit#(3))'(3'h1)));
                                writeLine_001 <= x_16;
                                victims_001 <= update (x_3, (Bit#(3))'(3'h5),
                                Struct25 {victim_valid : x_4, victim_idx :
                                (Bit#(3))'(3'h5), victim_line : x_16});

                            end else begin

                                Struct25 x_17 = ((x_3)[(Bit#(3))'(3'h6)]);
                                if (((x_17).victim_valid) &&
                                ((((x_17).victim_line).addr) ==
                                ((x_0).addr))) begin

                                    Struct24 x_18 = (Struct24 {addr :
                                    (x_0).addr, info_hit : (Bool)'(False),
                                    info_way : (x_0).info_way, info_write :
                                    (x_0).info_write, info : (x_0).info,
                                    value_write : (x_0).value_write, value :
                                    (x_0).value});
                                    writeStage_001 <= (x_4 ?
                                    ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h1)));

                                    writeLine_001 <= x_18;
                                    victims_001 <= update (x_3,
                                    (Bit#(3))'(3'h6), Struct25 {victim_valid
                                    : x_4, victim_idx : (Bit#(3))'(3'h6),
                                    victim_line : x_18});

                                end else begin

                                    Struct25 x_19 = ((x_3)[(Bit#(3))'(3'h7)]);

                                    if (((x_19).victim_valid) &&
                                    ((((x_19).victim_line).addr) ==
                                    ((x_0).addr))) begin

                                        Struct24 x_20 = (Struct24 {addr :
                                        (x_0).addr, info_hit :
                                        (Bool)'(False), info_way :
                                        (x_0).info_way, info_write :
                                        (x_0).info_write, info : (x_0).info,
                                        value_write : (x_0).value_write,
                                        value : (x_0).value});
                                        writeStage_001 <= (x_4 ?
                                        ((Bit#(3))'(3'h7)) :
                                        ((Bit#(3))'(3'h1)));
                                        writeLine_001 <= x_20;
                                        victims_001 <= update (x_3,
                                        (Bit#(3))'(3'h7), Struct25
                                        {victim_valid : x_4, victim_idx :
                                        (Bit#(3))'(3'h7), victim_line :
                                        x_20});

                                    end else begin

                                        writeStage_001 <= (Bit#(3))'(3'h1);

                                        writeLine_001 <= x_0;

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_001_writeRs ();
        let x_1 = (writeStage_001);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_001 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_001);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_001_hasVictimSlot ();
        let x_1 = (victims_001);
        Bool x_2 = ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) ||
        (((x_1)[(Bit#(3))'(3'h0)]).victim_valid))))))));
        return x_2;
    endmethod

    method ActionValue#(Struct24) cache_001_getVictim ();
        let x_1 = (victims_001);
        when ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid) ||
        (((x_1)[(Bit#(3))'(3'h0)]).victim_valid))))))), noAction);
        Struct24 x_2 = ((((x_1)[(Bit#(3))'(3'h7)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h7)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h6)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h6)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h5)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h5)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h4)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h4)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h3)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h3)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h2)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h2)]).victim_line) :
        ((((x_1)[(Bit#(3))'(3'h1)]).victim_valid ?
        (((x_1)[(Bit#(3))'(3'h1)]).victim_line) :
        (((x_1)[(Bit#(3))'(3'h0)]).victim_line)))))))))))))));
        return x_2;
    endmethod

    method Action cache_001_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_001);
        Struct25 x_2 = ((x_1)[(Bit#(3))'(3'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_001 <= update (x_1, (Bit#(3))'(3'h0),
            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct25 x_3 = ((x_1)[(Bit#(3))'(3'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_001 <= update (x_1, (Bit#(3))'(3'h1),
                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct25 x_4 = ((x_1)[(Bit#(3))'(3'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_001 <= update (x_1, (Bit#(3))'(3'h2),
                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct25 x_5 = ((x_1)[(Bit#(3))'(3'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_001 <= update (x_1, (Bit#(3))'(3'h3),
                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                        Struct25 x_6 = ((x_1)[(Bit#(3))'(3'h4)]);
                        if (((x_6).victim_valid) &&
                        ((((x_6).victim_line).addr) == (x_0))) begin

                            victims_001 <= update (x_1, (Bit#(3))'(3'h4),
                            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                        end else begin

                            Struct25 x_7 = ((x_1)[(Bit#(3))'(3'h5)]);
                            if (((x_7).victim_valid) &&
                            ((((x_7).victim_line).addr) == (x_0))) begin

                                victims_001 <= update (x_1, (Bit#(3))'(3'h5),
                                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                            end else begin

                                Struct25 x_8 = ((x_1)[(Bit#(3))'(3'h6)]);
                                if (((x_8).victim_valid) &&
                                ((((x_8).victim_line).addr) == (x_0))) begin

                                    victims_001 <= update (x_1,
                                    (Bit#(3))'(3'h6),
                                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                                end else begin

                                    Struct25 x_9 = ((x_1)[(Bit#(3))'(3'h7)]);

                                    if (((x_9).victim_valid) &&
                                    ((((x_9).victim_line).addr) == (x_0)))
                                    begin

                                        victims_001 <= update (x_1,
                                        (Bit#(3))'(3'h7),
                                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 3'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                                    end else begin

                                    end

                                end

                            end

                        end

                    end

                end

            end

        end

    endmethod

endmodule

interface Module146;
    method Action makeEnq_parentChildren001 (Struct10 x_0);
    method Action broadcast_parentChildren001 (Struct13 x_0);

endinterface


module mkModule146#(function Action enq_fifo00102(Struct2 _),
  function Action enq_fifo00112(Struct2 _),
  function Action enq_fifo00122(Struct2 _),
  function Action enq_fifo00132(Struct2 _),
  function Action enq_fifo0011(Struct2 _),
  function Action enq_fifo0010(Struct2 _)) (Module146);

    // No rules in this module

    method Action makeEnq_parentChildren001 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo0010((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo0011((x_0).enq_msg);

            end else begin

                Bit#(2) x_3 = ((x_0).enq_ch_idx);
                Struct2 x_4 = ((x_0).enq_msg);
                if ((x_3) == ((Bit#(2))'(2'h3))) begin
                let x_5 <- enq_fifo00132(x_4);

                end else begin

                    if ((x_3) == ((Bit#(2))'(2'h2))) begin
                    let x_6 <- enq_fifo00122(x_4);

                    end else begin

                        if ((x_3) == ((Bit#(2))'(2'h1))) begin
                        let x_7 <- enq_fifo00112(x_4);

                        end else begin

                            if ((x_3) == ((Bit#(2))'(2'h0))) begin
                            let x_8 <- enq_fifo00102(x_4);

                            end else begin

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method Action broadcast_parentChildren001 (Struct13 x_0);
        Bit#(4) x_1 = ((x_0).cs_inds);
        Struct2 x_2 = ((x_0).cs_msg);
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == (x_1))
        begin
        let x_3 <- enq_fifo00132(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == (x_1))
        begin
        let x_5 <- enq_fifo00122(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == (x_1))
        begin
        let x_7 <- enq_fifo00112(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == (x_1))
        begin
        let x_9 <- enq_fifo00102(x_2);

        end else begin

        end

    endmethod

endmodule

interface Module147;
    method Action cache_0010_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0010_readRs ();
    method Action cache_0010_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0010_writeRs ();
    method ActionValue#(Bool) cache_0010_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0010_getVictim ();
    method Action cache_0010_removeVictim (Bit#(64) x_0);

endinterface


module mkModule147#(function Action putRq_infoRam_0010_3(Struct36 _),
  function Action putRq_infoRam_0010_2(Struct36 _),
  function Action putRq_infoRam_0010_1(Struct36 _),
  function Action putRq_infoRam_0010_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0010(),
  function Action putRq_dataRam_0010(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0010_3(),
  function ActionValue#(Struct33) getRs_infoRam_0010_2(),
  function ActionValue#(Struct33) getRs_infoRam_0010_1(),
  function ActionValue#(Struct33) getRs_infoRam_0010_0()) (Module147);
    Reg#(Bit#(2)) readStage_0010 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0010 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0010 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0010 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0010 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0010 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0010 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0010 <- mkReg(unpack(0));

    rule read_tagmatch_0010;
        let x_0 = (readStage_0010);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0010);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0010_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0010_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0010_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0010_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0010 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0010 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0010(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0010 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0010;
        let x_0 = (readStage_0010);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0010 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0010();
        let x_2 = (readLine_0010);
        readLine_0010 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0010;
        let x_0 = (writeStage_0010);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0010);
        when ((x_1).info_hit, noAction);
        writeStage_0010 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0010_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0010_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0010_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0010_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0010(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0010;
        let x_0 = (writeStage_0010);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0010);
        when (! ((x_1).info_hit), noAction);
        writeStage_0010 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0010_0(x_4);
        let x_6 <- putRq_infoRam_0010_1(x_4);
        let x_7 <- putRq_infoRam_0010_2(x_4);
        let x_8 <- putRq_infoRam_0010_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0010;
        let x_0 = (writeStage_0010);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0010 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0010_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0010_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0010_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0010_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0010);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0010 <= x_10;
        victimLine_0010 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0010(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0010;
        let x_0 = (writeStage_0010);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0010);
        writeStage_0010 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0010);
        let x_6 = (victims_0010);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0010();
        let x_9 = (victimLine_0010);
        victims_0010 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0010 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0010_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0010_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0010_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0010_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0010(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0010_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0010);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0010);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0010);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0010 <= (Bit#(2))'(2'h3);
            readLine_0010 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0010 <= (Bit#(2))'(2'h3);
                readLine_0010 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0010 <= (Bit#(2))'(2'h3);
                    readLine_0010 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0010 <= (Bit#(2))'(2'h3);
                        readLine_0010 <= (x_7).victim_line;

                    end else begin

                        readStage_0010 <= (Bit#(2))'(2'h1);
                        readAddr_0010 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0010_0(x_9);
                        let x_11 <- putRq_infoRam_0010_1(x_9);
                        let x_12 <- putRq_infoRam_0010_2(x_9);
                        let x_13 <- putRq_infoRam_0010_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0010_readRs ();
        let x_1 = (readStage_0010);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0010 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0010);
        return x_2;
    endmethod

    method Action cache_0010_writeRq (Struct31 x_0);
        let x_1 = (readStage_0010);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0010);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0010);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0010 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0010 <= x_6;
            victims_0010 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0010 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0010 <= x_8;
                victims_0010 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0010 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0010 <= x_10;
                    victims_0010 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0010 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0010 <= x_12;
                        victims_0010 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0010 <= (Bit#(3))'(3'h1);
                        writeLine_0010 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0010_writeRs ();
        let x_1 = (writeStage_0010);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0010 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0010);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0010_hasVictimSlot ();
        let x_1 = (victims_0010);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0010_getVictim ();
        let x_1 = (victims_0010);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0010_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0010);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0010 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0010 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0010 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0010 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module148; method Action makeEnq_parentChildren0010 (Struct10 x_0);

endinterface


module mkModule148#(function Action enq_fifo001002(Struct2 _),
  function Action enq_fifo00101(Struct2 _),
  function Action enq_fifo00100(Struct2 _)) (Module148);

    // No rules in this module

    method Action makeEnq_parentChildren0010 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00100((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00101((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo001002(x_3);

            end

        end

    endmethod

endmodule

interface Module149;
    method Action cache_0011_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0011_readRs ();
    method Action cache_0011_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0011_writeRs ();
    method ActionValue#(Bool) cache_0011_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0011_getVictim ();
    method Action cache_0011_removeVictim (Bit#(64) x_0);

endinterface


module mkModule149#(function Action putRq_infoRam_0011_3(Struct36 _),
  function Action putRq_infoRam_0011_2(Struct36 _),
  function Action putRq_infoRam_0011_1(Struct36 _),
  function Action putRq_infoRam_0011_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0011(),
  function Action putRq_dataRam_0011(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0011_3(),
  function ActionValue#(Struct33) getRs_infoRam_0011_2(),
  function ActionValue#(Struct33) getRs_infoRam_0011_1(),
  function ActionValue#(Struct33) getRs_infoRam_0011_0()) (Module149);
    Reg#(Bit#(2)) readStage_0011 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0011 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0011 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0011 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0011 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0011 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0011 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0011 <- mkReg(unpack(0));

    rule read_tagmatch_0011;
        let x_0 = (readStage_0011);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0011);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0011_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0011_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0011_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0011_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0011 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0011 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0011(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0011 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0011;
        let x_0 = (readStage_0011);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0011 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0011();
        let x_2 = (readLine_0011);
        readLine_0011 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0011;
        let x_0 = (writeStage_0011);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0011);
        when ((x_1).info_hit, noAction);
        writeStage_0011 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0011_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0011_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0011_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0011_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0011(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0011;
        let x_0 = (writeStage_0011);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0011);
        when (! ((x_1).info_hit), noAction);
        writeStage_0011 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0011_0(x_4);
        let x_6 <- putRq_infoRam_0011_1(x_4);
        let x_7 <- putRq_infoRam_0011_2(x_4);
        let x_8 <- putRq_infoRam_0011_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0011;
        let x_0 = (writeStage_0011);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0011 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0011_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0011_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0011_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0011_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0011);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0011 <= x_10;
        victimLine_0011 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0011(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0011;
        let x_0 = (writeStage_0011);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0011);
        writeStage_0011 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0011);
        let x_6 = (victims_0011);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0011();
        let x_9 = (victimLine_0011);
        victims_0011 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0011 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0011_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0011_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0011_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0011_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0011(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0011_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0011);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0011);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0011);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0011 <= (Bit#(2))'(2'h3);
            readLine_0011 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0011 <= (Bit#(2))'(2'h3);
                readLine_0011 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0011 <= (Bit#(2))'(2'h3);
                    readLine_0011 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0011 <= (Bit#(2))'(2'h3);
                        readLine_0011 <= (x_7).victim_line;

                    end else begin

                        readStage_0011 <= (Bit#(2))'(2'h1);
                        readAddr_0011 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0011_0(x_9);
                        let x_11 <- putRq_infoRam_0011_1(x_9);
                        let x_12 <- putRq_infoRam_0011_2(x_9);
                        let x_13 <- putRq_infoRam_0011_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0011_readRs ();
        let x_1 = (readStage_0011);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0011 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0011);
        return x_2;
    endmethod

    method Action cache_0011_writeRq (Struct31 x_0);
        let x_1 = (readStage_0011);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0011);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0011);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0011 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0011 <= x_6;
            victims_0011 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0011 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0011 <= x_8;
                victims_0011 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0011 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0011 <= x_10;
                    victims_0011 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0011 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0011 <= x_12;
                        victims_0011 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0011 <= (Bit#(3))'(3'h1);
                        writeLine_0011 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0011_writeRs ();
        let x_1 = (writeStage_0011);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0011 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0011);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0011_hasVictimSlot ();
        let x_1 = (victims_0011);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0011_getVictim ();
        let x_1 = (victims_0011);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0011_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0011);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0011 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0011 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0011 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0011 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module150; method Action makeEnq_parentChildren0011 (Struct10 x_0);

endinterface


module mkModule150#(function Action enq_fifo001102(Struct2 _),
  function Action enq_fifo00111(Struct2 _),
  function Action enq_fifo00110(Struct2 _)) (Module150);

    // No rules in this module

    method Action makeEnq_parentChildren0011 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00110((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00111((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo001102(x_3);

            end

        end

    endmethod

endmodule

interface Module151;
    method Action cache_0012_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0012_readRs ();
    method Action cache_0012_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0012_writeRs ();
    method ActionValue#(Bool) cache_0012_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0012_getVictim ();
    method Action cache_0012_removeVictim (Bit#(64) x_0);

endinterface


module mkModule151#(function Action putRq_infoRam_0012_3(Struct36 _),
  function Action putRq_infoRam_0012_2(Struct36 _),
  function Action putRq_infoRam_0012_1(Struct36 _),
  function Action putRq_infoRam_0012_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0012(),
  function Action putRq_dataRam_0012(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0012_3(),
  function ActionValue#(Struct33) getRs_infoRam_0012_2(),
  function ActionValue#(Struct33) getRs_infoRam_0012_1(),
  function ActionValue#(Struct33) getRs_infoRam_0012_0()) (Module151);
    Reg#(Bit#(2)) readStage_0012 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0012 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0012 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0012 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0012 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0012 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0012 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0012 <- mkReg(unpack(0));

    rule read_tagmatch_0012;
        let x_0 = (readStage_0012);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0012);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0012_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0012_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0012_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0012_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0012 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0012 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0012(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0012 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0012;
        let x_0 = (readStage_0012);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0012 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0012();
        let x_2 = (readLine_0012);
        readLine_0012 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0012;
        let x_0 = (writeStage_0012);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0012);
        when ((x_1).info_hit, noAction);
        writeStage_0012 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0012_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0012_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0012_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0012_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0012(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0012;
        let x_0 = (writeStage_0012);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0012);
        when (! ((x_1).info_hit), noAction);
        writeStage_0012 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0012_0(x_4);
        let x_6 <- putRq_infoRam_0012_1(x_4);
        let x_7 <- putRq_infoRam_0012_2(x_4);
        let x_8 <- putRq_infoRam_0012_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0012;
        let x_0 = (writeStage_0012);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0012 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0012_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0012_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0012_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0012_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0012);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0012 <= x_10;
        victimLine_0012 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0012(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0012;
        let x_0 = (writeStage_0012);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0012);
        writeStage_0012 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0012);
        let x_6 = (victims_0012);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0012();
        let x_9 = (victimLine_0012);
        victims_0012 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0012 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0012_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0012_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0012_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0012_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0012(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0012_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0012);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0012);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0012);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0012 <= (Bit#(2))'(2'h3);
            readLine_0012 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0012 <= (Bit#(2))'(2'h3);
                readLine_0012 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0012 <= (Bit#(2))'(2'h3);
                    readLine_0012 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0012 <= (Bit#(2))'(2'h3);
                        readLine_0012 <= (x_7).victim_line;

                    end else begin

                        readStage_0012 <= (Bit#(2))'(2'h1);
                        readAddr_0012 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0012_0(x_9);
                        let x_11 <- putRq_infoRam_0012_1(x_9);
                        let x_12 <- putRq_infoRam_0012_2(x_9);
                        let x_13 <- putRq_infoRam_0012_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0012_readRs ();
        let x_1 = (readStage_0012);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0012 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0012);
        return x_2;
    endmethod

    method Action cache_0012_writeRq (Struct31 x_0);
        let x_1 = (readStage_0012);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0012);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0012);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0012 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0012 <= x_6;
            victims_0012 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0012 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0012 <= x_8;
                victims_0012 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0012 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0012 <= x_10;
                    victims_0012 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0012 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0012 <= x_12;
                        victims_0012 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0012 <= (Bit#(3))'(3'h1);
                        writeLine_0012 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0012_writeRs ();
        let x_1 = (writeStage_0012);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0012 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0012);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0012_hasVictimSlot ();
        let x_1 = (victims_0012);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0012_getVictim ();
        let x_1 = (victims_0012);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0012_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0012);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0012 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0012 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0012 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0012 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module152; method Action makeEnq_parentChildren0012 (Struct10 x_0);

endinterface


module mkModule152#(function Action enq_fifo001202(Struct2 _),
  function Action enq_fifo00121(Struct2 _),
  function Action enq_fifo00120(Struct2 _)) (Module152);

    // No rules in this module

    method Action makeEnq_parentChildren0012 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00120((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00121((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo001202(x_3);

            end

        end

    endmethod

endmodule

interface Module153;
    method Action cache_0013_readRq (Bit#(64) x_0);
    method ActionValue#(Struct31) cache_0013_readRs ();
    method Action cache_0013_writeRq (Struct31 x_0);
    method ActionValue#(Struct31) cache_0013_writeRs ();
    method ActionValue#(Bool) cache_0013_hasVictimSlot ();
    method ActionValue#(Struct31) cache_0013_getVictim ();
    method Action cache_0013_removeVictim (Bit#(64) x_0);

endinterface


module mkModule153#(function Action putRq_infoRam_0013_3(Struct36 _),
  function Action putRq_infoRam_0013_2(Struct36 _),
  function Action putRq_infoRam_0013_1(Struct36 _),
  function Action putRq_infoRam_0013_0(Struct36 _),
  function ActionValue#(Bit#(64)) getRs_dataRam_0013(),
  function Action putRq_dataRam_0013(Struct35 _),
  function ActionValue#(Struct33) getRs_infoRam_0013_3(),
  function ActionValue#(Struct33) getRs_infoRam_0013_2(),
  function ActionValue#(Struct33) getRs_infoRam_0013_1(),
  function ActionValue#(Struct33) getRs_infoRam_0013_0()) (Module153);
    Reg#(Bit#(2)) readStage_0013 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_0013 <- mkReg(unpack(0));
    Reg#(Struct31) readLine_0013 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_0013 <- mkReg(unpack(0));
    Reg#(Struct31) writeLine_0013 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct32)) victims_0013 <- mkReg(unpack(0));
    Reg#(Struct31) victimLine_0013 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_0013 <- mkReg(unpack(0));

    rule read_tagmatch_0013;
        let x_0 = (readStage_0013);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_0013);
        Bit#(55) x_2 = ((x_1)[63:9]);
        Bit#(6) x_3 = ((x_1)[8:3]);
        Vector#(4, Struct33) x_4 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_0013_0();
        Vector#(4, Struct33) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_0013_1();
        Vector#(4, Struct33) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_0013_2();
        Vector#(4, Struct33) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_0013_3();
        Vector#(4, Struct33) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct34 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct34 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct34 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct34)'(Struct34 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_0013 <= Struct31 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Bit#(64))'(64'h0)};
        if ((x_13).tm_hit) begin

            readStage_0013 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_0013(Struct35 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain : (Bit#(64))'(64'h0)});

        end else begin
        readStage_0013 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_0013;
        let x_0 = (readStage_0013);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_0013 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_0013();
        let x_2 = (readLine_0013);
        readLine_0013 <= Struct31 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_0013;
        let x_0 = (writeStage_0013);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0013);
        when ((x_1).info_hit, noAction);
        writeStage_0013 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct36 x_6 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_0013_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_0013_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_0013_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_0013_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_0013(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_0013;
        let x_0 = (writeStage_0013);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_0013);
        when (! ((x_1).info_hit), noAction);
        writeStage_0013 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(6) x_3 = ((x_2)[8:3]);
        Struct36 x_4 = (Struct36 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_0013_0(x_4);
        let x_6 <- putRq_infoRam_0013_1(x_4);
        let x_7 <- putRq_infoRam_0013_2(x_4);
        let x_8 <- putRq_infoRam_0013_3(x_4);

    endrule

    rule write_info_miss_rep_rs_0013;
        let x_0 = (writeStage_0013);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_0013 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct33) x_1 =
        ((Vector#(4, Struct33))'(vec(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_0013_0();
        Vector#(4, Struct33) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_0013_1();
        Vector#(4, Struct33) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_0013_2();
        Vector#(4, Struct33) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_0013_3();
        Vector#(4, Struct33) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_0013);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(6) x_13 = ((x_12)[8:3]);
        Struct33 x_14 = ((x_9)[x_10]);
        Bit#(55) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_0013 <= x_10;
        victimLine_0013 <= Struct31 {addr :
        {(x_15),({(x_13),((Bit#(3))'(3'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value : (Bit#(64))'(64'h0)};
        let x_17 <- putRq_dataRam_0013(Struct35 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain : (Bit#(64))'(64'h0)});

    endrule

    rule write_victim_rs_0013;
        let x_0 = (writeStage_0013);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_0013);
        writeStage_0013 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(55) x_3 = ((x_2)[63:9]);
        Bit#(6) x_4 = ((x_2)[8:3]);
        let x_5 = (victimWay_0013);
        let x_6 = (victims_0013);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_0013();
        let x_9 = (victimLine_0013);
        victims_0013 <= update (x_6, x_7, Struct32 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct31 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_0013 <= Struct31 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct36 x_10 = (Struct36 {write : (Bool)'(True), addr : x_4,
            datain : Struct33 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_0013_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_0013_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_0013_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_0013_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_0013(Struct35 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_0013_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_0013);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_0013);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_0013);
        Struct32 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin

            readStage_0013 <= (Bit#(2))'(2'h3);
            readLine_0013 <= (x_4).victim_line;

        end else begin

            Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_0013 <= (Bit#(2))'(2'h3);
                readLine_0013 <= (x_5).victim_line;

            end else begin

                Struct32 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_0013 <= (Bit#(2))'(2'h3);
                    readLine_0013 <= (x_6).victim_line;

                end else begin

                    Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_0013 <= (Bit#(2))'(2'h3);
                        readLine_0013 <= (x_7).victim_line;

                    end else begin

                        readStage_0013 <= (Bit#(2))'(2'h1);
                        readAddr_0013 <= x_0;
                        Bit#(6) x_8 = ((x_0)[8:3]);
                        Struct36 x_9 = (Struct36 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct33)'(Struct33 {tag: 55'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_0013_0(x_9);
                        let x_11 <- putRq_infoRam_0013_1(x_9);
                        let x_12 <- putRq_infoRam_0013_2(x_9);
                        let x_13 <- putRq_infoRam_0013_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0013_readRs ();
        let x_1 = (readStage_0013);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_0013 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_0013);
        return x_2;
    endmethod

    method Action cache_0013_writeRq (Struct31 x_0);
        let x_1 = (readStage_0013);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_0013);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_0013);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct32 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct31 x_6 = (Struct31 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_0013 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_0013 <= x_6;
            victims_0013 <= update (x_3, (Bit#(2))'(2'h0), Struct32
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct32 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct31 x_8 = (Struct31 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_0013 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_0013 <= x_8;
                victims_0013 <= update (x_3, (Bit#(2))'(2'h1), Struct32
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct32 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct31 x_10 = (Struct31 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_0013 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_0013 <= x_10;
                    victims_0013 <= update (x_3, (Bit#(2))'(2'h2), Struct32
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct32 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct31 x_12 = (Struct31 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_0013 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_0013 <= x_12;
                        victims_0013 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct32 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin

                        writeStage_0013 <= (Bit#(3))'(3'h1);
                        writeLine_0013 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct31) cache_0013_writeRs ();
        let x_1 = (writeStage_0013);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_0013 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_0013);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_0013_hasVictimSlot ();
        let x_1 = (victims_0013);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct31) cache_0013_getVictim ();
        let x_1 = (victims_0013);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct31 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_0013_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_0013);
        Struct32 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_0013 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


        end else begin

            Struct32 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_0013 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


            end else begin

                Struct32 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_0013 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                end else begin

                    Struct32 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_0013 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct32)'(Struct32 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module154; method Action makeEnq_parentChildren0013 (Struct10 x_0);

endinterface


module mkModule154#(function Action enq_fifo001302(Struct2 _),
  function Action enq_fifo00131(Struct2 _),
  function Action enq_fifo00130(Struct2 _)) (Module154);

    // No rules in this module

    method Action makeEnq_parentChildren0013 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo00130((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo00131((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo001302(x_3);

            end

        end

    endmethod

endmodule

interface Module155;
endinterface


module mkModule155#(function ActionValue#(Struct3) cache_00_writeRs(),
  function Action cache_00_removeVictim(Bit#(64) _),
  function ActionValue#(Struct3) cache_00_getVictim(),
  function Action transferUpDown00(Struct17 _),
  function Action releaseDL00(Bit#(64) _),
  function Action releaseUL00(Bit#(64) _),
  function ActionValue#(Struct15) upLockGet00(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0011(),
  function Action addRs00(Struct14 _),
  function ActionValue#(Struct6) downLockGet00(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0001(),
  function Action broadcast_parentChildren00(Struct13 _),
  function Action registerDL00(Struct12 _),
  function Action registerUL00(Struct11 _),
  function ActionValue#(Bool) cache_00_hasVictimSlot(),
  function Action makeEnq_parentChildren00(Struct10 _),
  function Action cache_00_writeRq(Struct3 _),
  function ActionValue#(Bool) downLockable00(Bit#(64) _),
  function ActionValue#(Bool) upLockable00(Bit#(64) _),
  function ActionValue#(Struct3) cache_00_readRs(),
  function ActionValue#(Struct2) deq_fifo0010(),
  function ActionValue#(Struct2) deq_fifo0000(),
  function ActionValue#(Struct6) downLockRssFull00(),
  function Action cache_00_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo002()) (Module155);
    Reg#(Bit#(2)) rr00 <- mkReg(unpack(0));
    Reg#(Struct1) prl00 <- mkReg(unpack(0));
    Reg#(Struct1) crqrl00 <- mkReg(unpack(0));
    Reg#(Struct1) crsrl00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc00 <- mkReg(unpack(0));
    Reg#(Struct5) wl00 <- mkReg(unpack(0));

    rule rr_00;let x_0 = (rr00);
               rr00 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_00_1230;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo002();
        prl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc00 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_1232;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull00();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc00 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_00_readRq((x_4).addr);

    endrule

    rule rule_00_12310000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo0000();
        crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc00 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_12310010;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo0010();
        crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h1), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc00 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_456;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        let x_3 <- cache_00_readRs();
        let x_4 = (rlc00);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl00 <= Struct1 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl00 <= Struct1 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl00 <= Struct1 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_00_000000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_001000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_01000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_03000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_10000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 = (wl00);
        when (! ((x_23).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_14000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_15000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))), r_dl_rsbTo : (Bit#(4))'(4'h8)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_25000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_2600000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_2601000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_261000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_27000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_28000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_290000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_291000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_210000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_211000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_00_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_040000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_070000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1600000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1601000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11000000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11001000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11002000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_000001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_001001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_01001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_03001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_10001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 = (wl00);
        when (! ((x_23).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_14001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_15001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))), r_dl_rsbTo : (Bit#(4))'(4'h9)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_25001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_2600001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_2601001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_261001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_27001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_28001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_290001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_291001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_210001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_211001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_00_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_040001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_070001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1600001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1601001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11000001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11001001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11002001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        Struct3 x_4 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo0011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet00((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs00(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_020;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_19 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct3 x_22 = (Struct3 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_00_writeRq(x_22);
        let x_24 <- releaseUL00((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren00(x_25);
        let x_27 = (wl00);
        when (! ((x_27).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_021;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_19 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct3 x_22 = (Struct3 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_00_writeRq(x_22);
        let x_24 <- releaseUL00((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren00(x_25);
        let x_27 = (wl00);
        when (! ((x_27).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_041;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct3 x_18 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_st,
        mesi_dir_sharers : (((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_sharers) :
        (((Bit#(4))'(4'h1)) << ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_00_writeRq(x_21);
        let x_23 <- releaseDL00((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 = (wl00);
        when (! ((x_26).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_05;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_10).dir_st))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct3 x_16 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_17 = (Struct3 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_06;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_9))) && ((!
        (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_10).dir_st))))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_071;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct3 x_18 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0),
        dir_sharers : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (x_20).info_write, info : (x_20).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        let x_22 <- cache_00_writeRq(x_21);
        let x_23 <- releaseDL00((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 = (wl00);
        when (! ((x_26).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_12;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((x_10).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))), noAction);

        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_19 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_00_writeRq(x_21);
        let x_23 <- releaseUL00((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 = (wl00);
        when (! ((x_26).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_13;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))) ==
        ((Bit#(4))'(4'h0)))) && (((x_10).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = ((x_13).ul_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_18 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_19 <- cache_00_writeRq(x_18);
        let x_20 <- transferUpDown00(Struct17 {r_dl_addr : (x_11).addr,
        r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))});
        let x_21 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((x_17)[1:0]))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_16).addr, value : (Bit#(64))'(64'h0)}});
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_161;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        let x_21 <- releaseDL00((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_170;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_10).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct3 x_16 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_17 = (Struct3 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_171;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct3 x_16 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_17 = (Struct3 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_190;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_191;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_192;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11010;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        let x_21 <- releaseDL00((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11011;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        let x_21 <- releaseDL00((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_20;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        let x_4 <- cache_00_getVictim();
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_9))
        && ((x_9) < ((Bit#(3))'(3'h4)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        let x_15 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren00(x_16);
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_21;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        let x_4 <- cache_00_getVictim();
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when ((((x_10).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_8) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_9))) || (((x_8) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) && ((x_9) <
        ((Bit#(3))'(3'h3)))))), noAction);
        let x_15 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren00(x_16);
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_22;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL00((x_11).addr);
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_00_removeVictim(x_19);
        let x_21 = (crqrl00);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl00 <= Struct1 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct3 {addr : x_19, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl00);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl00 <= Struct1 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct3 {addr : x_19, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    (* descending_urgency = "rule_00_23, rule_00_20, rule_00_21" *)
    rule rule_00_23;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        let x_4 <- cache_00_getVictim();
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((x_9) == ((Bit#(3))'(3'h1))) && (! (((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_9) == ((Bit#(3))'(3'h2))) && ((x_8) ==
        ((Bool)'(False)))), noAction);
        let x_16 = (wl00);
        when (! ((x_16).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_17 = ((x_11).addr);
        let x_18 <- cache_00_removeVictim(x_17);
        let x_19 = (crqrl00);
        if ((((x_19).rl_valid) && ((x_19).rl_line_valid)) &&
        ((((x_19).rl_msg).addr) == (x_17))) begin

            crqrl00 <= Struct1 {rl_valid : (x_19).rl_valid, rl_cmidx :
            (x_19).rl_cmidx, rl_msg : (x_19).rl_msg, rl_line_valid :
            (x_19).rl_line_valid, rl_line : Struct3 {addr : x_17, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_21 = (crsrl00);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_17))) begin

            crsrl00 <= Struct1 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct3 {addr : x_17, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_00_7890;
        let x_0 = (wl00);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl00 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_00_7891;
        let x_0 = (wl00);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_00_writeRs();
        let x_2 = (prl00);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl00);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl00);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl00 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module156;
endinterface


module mkModule156#(function ActionValue#(Struct24) cache_000_writeRs(),
  function Action cache_000_removeVictim(Bit#(64) _),
  function ActionValue#(Struct24) cache_000_getVictim(),
  function Action transferUpDown000(Struct17 _),
  function Action releaseDL000(Bit#(64) _),
  function Action releaseUL000(Bit#(64) _),
  function ActionValue#(Struct15) upLockGet000(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00031(),
  function ActionValue#(Struct2) deq_fifo00021(),
  function ActionValue#(Struct2) deq_fifo00011(),
  function Action addRs000(Struct14 _),
  function ActionValue#(Struct6) downLockGet000(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00001(),
  function Action broadcast_parentChildren000(Struct13 _),
  function Action registerDL000(Struct12 _),
  function Action registerUL000(Struct11 _),
  function ActionValue#(Bool) cache_000_hasVictimSlot(),
  function Action makeEnq_parentChildren000(Struct10 _),
  function Action cache_000_writeRq(Struct24 _),
  function ActionValue#(Bool) downLockable000(Bit#(64) _),
  function ActionValue#(Bool) upLockable000(Bit#(64) _),
  function ActionValue#(Struct24) cache_000_readRs(),
  function ActionValue#(Struct2) deq_fifo00030(),
  function ActionValue#(Struct2) deq_fifo00020(),
  function ActionValue#(Struct2) deq_fifo00010(),
  function ActionValue#(Struct2) deq_fifo00000(),
  function ActionValue#(Struct6) downLockRssFull000(),
  function Action cache_000_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0002()) (Module156);
    Reg#(Bit#(2)) rr000 <- mkReg(unpack(0));
    Reg#(Struct23) prl000 <- mkReg(unpack(0));
    Reg#(Struct23) crqrl000 <- mkReg(unpack(0));
    Reg#(Struct23) crsrl000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc000 <- mkReg(unpack(0));
    Reg#(Struct5) wl000 <- mkReg(unpack(0));

    rule rr_000;let x_0 = (rr000);
                rr000 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_000_1230;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo0002();
        prl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc000 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_000_readRq((x_3).addr);

    endrule

    rule rule_000_1232;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull000();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc000 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_000_readRq((x_4).addr);

    endrule

    rule rule_000_123100000;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00000();
        crqrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc000 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_000_readRq((x_3).addr);

    endrule

    rule rule_000_123100010;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00010();
        crqrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h1), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc000 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_000_readRq((x_3).addr);

    endrule

    rule rule_000_123100020;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00020();
        crqrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h2), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc000 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_000_readRq((x_3).addr);

    endrule

    rule rule_000_123100030;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00030();
        crqrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h3), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc000 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_000_readRq((x_3).addr);

    endrule

    rule rule_000_456;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        let x_3 <- cache_000_readRs();
        let x_4 = (rlc000);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl000 <= Struct23 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl000 <= Struct23 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl000 <= Struct23 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_000_0000000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0010000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_010000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_030000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_100000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
        let x_23 = (wl000);
        when (! ((x_23).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_110000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_140000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_150000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        let x_17 <- broadcast_parentChildren000(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_250000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_26000000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_26010000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2610000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_270000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_280000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_2900000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2910000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2100000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2110000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_000_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 = (wl000);
        when (! ((x_24).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0400000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_0700000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16000000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16010000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110000000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110010000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110020000;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00001();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_0000001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0010001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_010001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_030001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_100001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
        let x_23 = (wl000);
        when (! ((x_23).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_110001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_140001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_150001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        let x_17 <- broadcast_parentChildren000(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_250001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_26000001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_26010001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2610001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_270001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_280001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_2900001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2910001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2100001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2110001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_000_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 = (wl000);
        when (! ((x_24).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0400001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_0700001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16000001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16010001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110000001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110010001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110020001;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00011();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_0000002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0010002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_010002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_030002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_100002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
        let x_23 = (wl000);
        when (! ((x_23).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_110002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_140002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_150002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        let x_17 <- broadcast_parentChildren000(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_250002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_26000002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_26010002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2610002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_270002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_280002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_2900002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2910002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2100002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2110002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_000_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 = (wl000);
        when (! ((x_24).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0400002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00021();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_0700002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00021();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16000002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00021();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16010002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00021();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110000002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00021();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110010002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00021();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110020002;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00021();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_0000003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0010003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_010003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_030003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_100003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren000(x_21);
        let x_23 = (wl000);
        when (! ((x_23).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_110003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_140003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_150003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        let x_17 <- broadcast_parentChildren000(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_250003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_26000003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_26010003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2610003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_270003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_280003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_2900003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2910003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2100003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_000_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren000(x_20);
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_2110003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_000_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 = (wl000);
        when (! ((x_24).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_0400003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00031();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_0700003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00031();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16000003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00031();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_16010003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00031();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110000003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00031();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110010003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00031();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_110020003;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00031();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet000((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs000(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_020;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct24 x_22 = (Struct24 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_000_writeRq(x_22);
        let x_24 <- releaseUL000((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren000(x_25);
        let x_27 = (wl000);
        when (! ((x_27).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_021;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct24 x_22 = (Struct24 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_000_writeRq(x_22);
        let x_24 <- releaseUL000((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren000(x_25);
        let x_27 = (wl000);
        when (! ((x_27).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_041;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet000((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct24 x_18 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_st,
        mesi_dir_sharers : (((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_sharers) :
        (((Bit#(4))'(4'h1)) << ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_000_writeRq(x_21);
        let x_23 <- releaseDL000((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren000(x_24);
        let x_26 = (wl000);
        when (! ((x_26).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_05;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_10).dir_st))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_06;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_9))) && ((!
        (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_10).dir_st))))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_071;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet000((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct24 x_18 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0),
        dir_sharers : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (x_20).info_write, info : (x_20).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        let x_22 <- cache_000_writeRq(x_21);
        let x_23 <- releaseDL000((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren000(x_24);
        let x_26 = (wl000);
        when (! ((x_26).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_12;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((x_10).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))), noAction);

        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_000_writeRq(x_21);
        let x_23 <- releaseUL000((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren000(x_24);
        let x_26 = (wl000);
        when (! ((x_26).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_13;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))) ==
        ((Bit#(4))'(4'h0)))) && (((x_10).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = ((x_13).ul_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_18 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_19 <- cache_000_writeRq(x_18);
        let x_20 <- transferUpDown000(Struct17 {r_dl_addr : (x_11).addr,
        r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))});
        let x_21 <- broadcast_parentChildren000(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((x_17)[1:0]))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_16).addr, value : (Bit#(64))'(64'h0)}});
        let x_22 = (wl000);
        when (! ((x_22).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_161;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet000((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        let x_21 <- releaseDL000((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 = (wl000);
        when (! ((x_24).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_170;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_10).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_171;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_190;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_17 <- broadcast_parentChildren000(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_191;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_192;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL000(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_17 <- broadcast_parentChildren000(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_11010;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet000((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        let x_21 <- releaseDL000((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 = (wl000);
        when (! ((x_24).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_11011;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet000((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        let x_21 <- releaseDL000((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren000(x_22);
        let x_24 = (wl000);
        when (! ((x_24).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_20;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        let x_4 <- cache_000_getVictim();
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_9))
        && ((x_9) < ((Bit#(3))'(3'h4)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        let x_15 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren000(x_16);
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_21;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        let x_4 <- cache_000_getVictim();
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when ((((x_10).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_8) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_9))) || (((x_8) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) && ((x_9) <
        ((Bit#(3))'(3'h3)))))), noAction);
        let x_15 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren000(x_16);
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_22;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL000((x_11).addr);
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_000_removeVictim(x_19);
        let x_21 = (crqrl000);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl000 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl000);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl000 <= Struct23 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    (* descending_urgency = "rule_000_23, rule_000_20, rule_000_21" *)
    rule rule_000_23;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        let x_4 <- cache_000_getVictim();
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((((x_9) == ((Bit#(3))'(3'h1))) && (! (((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_9) == ((Bit#(3))'(3'h2))) && ((x_8) ==
        ((Bool)'(False)))), noAction);
        let x_16 = (wl000);
        when (! ((x_16).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_17 = ((x_11).addr);
        let x_18 <- cache_000_removeVictim(x_17);
        let x_19 = (crqrl000);
        if ((((x_19).rl_valid) && ((x_19).rl_line_valid)) &&
        ((((x_19).rl_msg).addr) == (x_17))) begin

            crqrl000 <= Struct23 {rl_valid : (x_19).rl_valid, rl_cmidx :
            (x_19).rl_cmidx, rl_msg : (x_19).rl_msg, rl_line_valid :
            (x_19).rl_line_valid, rl_line : Struct24 {addr : x_17, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_21 = (crsrl000);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_17))) begin

            crsrl000 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_17, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_000_7890;
        let x_0 = (wl000);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl000 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_000_7891;
        let x_0 = (wl000);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_000_writeRs();
        let x_2 = (prl000);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl000);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl000);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl000 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module157;
endinterface


module mkModule157#(function ActionValue#(Struct31) cache_0000_writeRs(),
  function Action cache_0000_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0000_getVictim(),
  function Action releaseUL0000(Bit#(64) _),
  function Action cache_0000_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0000(Bit#(64) _),
  function Action registerUL0000(Struct11 _),
  function ActionValue#(Bool) cache_0000_hasVictimSlot(),
  function Action makeEnq_parentChildren0000(Struct10 _),
  function ActionValue#(Bool) downLockable0000(Bit#(64) _),
  function ActionValue#(Bool) upLockable0000(Bit#(64) _),
  function ActionValue#(Struct31) cache_0000_readRs(),
  function ActionValue#(Struct2) deq_fifo000000(),
  function ActionValue#(Struct6) downLockRssFull0000(),
  function Action cache_0000_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00002()) (Module157);
    Reg#(Bit#(2)) rr0000 <- mkReg(unpack(0));
    Reg#(Struct30) prl0000 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0000 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0000 <- mkReg(unpack(0));
    Reg#(Struct5) wl0000 <- mkReg(unpack(0));

    rule rr_0000;let x_0 = (rr0000);
                 rr0000 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0000_1230;
        let x_0 = (prl0000);
        let x_1 = (crqrl0000);
        let x_2 = (crsrl0000);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00002();
        prl0000 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0000 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0000_readRq((x_3).addr);

    endrule

    rule rule_0000_1232;
        let x_0 = (prl0000);
        let x_1 = (crqrl0000);
        let x_2 = (crsrl0000);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0000();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0000 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0000 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0000_readRq((x_4).addr);

    endrule

    rule rule_0000_1231000000;
        let x_0 = (prl0000);
        let x_1 = (crqrl0000);
        let x_2 = (crsrl0000);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo000000();
        crqrl0000 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0000 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0000_readRq((x_3).addr);

    endrule

    rule rule_0000_456;
        let x_0 = (prl0000);
        let x_1 = (crqrl0000);
        let x_2 = (crsrl0000);
        let x_3 <- cache_0000_readRs();
        let x_4 = (rlc0000);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0000 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0000 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0000 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0000_00;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0000((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0000(x_17);
        let x_19 = (wl0000);
        when (! ((x_19).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0000_01;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0000((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0000(x_18);
        let x_20 = (wl0000);
        when (! ((x_20).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0000_020;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0000_writeRq(x_20);
        let x_22 <- releaseUL0000((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0000(x_23);
        let x_25 = (wl0000);
        when (! ((x_25).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_021;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0000_writeRq(x_20);
        let x_22 <- releaseUL0000((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0000(x_23);
        let x_25 = (wl0000);
        when (! ((x_25).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_03;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0000((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0000(x_19);
        let x_21 = (wl0000);
        when (! ((x_21).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_100;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0000((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0000_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0000(x_21);
        let x_23 = (wl0000);
        when (! ((x_23).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_101;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0000(x_19);
        let x_21 = (wl0000);
        when (! ((x_21).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_11;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0000((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0000(x_18);
        let x_20 = (wl0000);
        when (! ((x_20).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0000_12;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0000_writeRq(x_21);
        let x_23 <- releaseUL0000((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0000(x_24);
        let x_26 = (wl0000);
        when (! ((x_26).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_130;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0000((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0000(x_19);
        let x_21 = (wl0000);
        when (! ((x_21).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_131;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0000((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0000(x_19);
        let x_21 = (wl0000);
        when (! ((x_21).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0000_20;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        let x_4 <- cache_0000_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0000((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0000(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0000(x_16);
        let x_18 = (wl0000);
        when (! ((x_18).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0000_20, rule_0000_21" *)
    rule rule_0000_21;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        let x_4 <- cache_0000_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0000((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0000(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0000(x_16);
        let x_18 = (wl0000);
        when (! ((x_18).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0000_22;
        let x_0 = (rr0000);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0000);
        let x_2 = (crqrl0000);
        let x_3 = (crsrl0000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0000 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0000((x_11).addr);
        let x_18 = (wl0000);
        when (! ((x_18).wl_valid), noAction);
        wl0000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0000_removeVictim(x_19);
        let x_21 = (crqrl0000);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0000 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0000);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0000 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0000_7890;
        let x_0 = (wl0000);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0000 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0000_7891;
        let x_0 = (wl0000);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0000_writeRs();
        let x_2 = (prl0000);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0000 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0000);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0000 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0000);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0000 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0000 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module158;
endinterface


module mkModule158#(function ActionValue#(Struct31) cache_0001_writeRs(),
  function Action cache_0001_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0001_getVictim(),
  function Action releaseUL0001(Bit#(64) _),
  function Action cache_0001_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0001(Bit#(64) _),
  function Action registerUL0001(Struct11 _),
  function ActionValue#(Bool) cache_0001_hasVictimSlot(),
  function Action makeEnq_parentChildren0001(Struct10 _),
  function ActionValue#(Bool) downLockable0001(Bit#(64) _),
  function ActionValue#(Bool) upLockable0001(Bit#(64) _),
  function ActionValue#(Struct31) cache_0001_readRs(),
  function ActionValue#(Struct2) deq_fifo000100(),
  function ActionValue#(Struct6) downLockRssFull0001(),
  function Action cache_0001_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00012()) (Module158);
    Reg#(Bit#(2)) rr0001 <- mkReg(unpack(0));
    Reg#(Struct30) prl0001 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0001 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0001 <- mkReg(unpack(0));
    Reg#(Struct5) wl0001 <- mkReg(unpack(0));

    rule rr_0001;let x_0 = (rr0001);
                 rr0001 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0001_1230;
        let x_0 = (prl0001);
        let x_1 = (crqrl0001);
        let x_2 = (crsrl0001);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00012();
        prl0001 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0001 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0001_readRq((x_3).addr);

    endrule

    rule rule_0001_1232;
        let x_0 = (prl0001);
        let x_1 = (crqrl0001);
        let x_2 = (crsrl0001);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0001();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0001 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0001 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0001_readRq((x_4).addr);

    endrule

    rule rule_0001_1231000100;
        let x_0 = (prl0001);
        let x_1 = (crqrl0001);
        let x_2 = (crsrl0001);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo000100();
        crqrl0001 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0001 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0001_readRq((x_3).addr);

    endrule

    rule rule_0001_456;
        let x_0 = (prl0001);
        let x_1 = (crqrl0001);
        let x_2 = (crsrl0001);
        let x_3 <- cache_0001_readRs();
        let x_4 = (rlc0001);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0001 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0001 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0001 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0001_00;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0001((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0001(x_17);
        let x_19 = (wl0001);
        when (! ((x_19).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0001_01;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0001((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0001(x_18);
        let x_20 = (wl0001);
        when (! ((x_20).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0001_020;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0001_writeRq(x_20);
        let x_22 <- releaseUL0001((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0001(x_23);
        let x_25 = (wl0001);
        when (! ((x_25).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_021;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0001_writeRq(x_20);
        let x_22 <- releaseUL0001((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0001(x_23);
        let x_25 = (wl0001);
        when (! ((x_25).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_03;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0001((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0001(x_19);
        let x_21 = (wl0001);
        when (! ((x_21).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_100;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0001((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0001_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0001(x_21);
        let x_23 = (wl0001);
        when (! ((x_23).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_101;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0001(x_19);
        let x_21 = (wl0001);
        when (! ((x_21).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_11;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0001((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0001(x_18);
        let x_20 = (wl0001);
        when (! ((x_20).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0001_12;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0001_writeRq(x_21);
        let x_23 <- releaseUL0001((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0001(x_24);
        let x_26 = (wl0001);
        when (! ((x_26).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_130;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0001((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0001(x_19);
        let x_21 = (wl0001);
        when (! ((x_21).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_131;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0001((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0001(x_19);
        let x_21 = (wl0001);
        when (! ((x_21).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0001_20;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        let x_4 <- cache_0001_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0001(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0001(x_16);
        let x_18 = (wl0001);
        when (! ((x_18).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0001_20, rule_0001_21" *)
    rule rule_0001_21;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        let x_4 <- cache_0001_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0001((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0001(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0001(x_16);
        let x_18 = (wl0001);
        when (! ((x_18).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0001_22;
        let x_0 = (rr0001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0001);
        let x_2 = (crqrl0001);
        let x_3 = (crsrl0001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0001 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0001((x_11).addr);
        let x_18 = (wl0001);
        when (! ((x_18).wl_valid), noAction);
        wl0001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0001_removeVictim(x_19);
        let x_21 = (crqrl0001);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0001 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0001);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0001 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0001_7890;
        let x_0 = (wl0001);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0001 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0001_7891;
        let x_0 = (wl0001);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0001_writeRs();
        let x_2 = (prl0001);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0001 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0001);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0001 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0001);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0001 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0001 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module159;
endinterface


module mkModule159#(function ActionValue#(Struct31) cache_0002_writeRs(),
  function Action cache_0002_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0002_getVictim(),
  function Action releaseUL0002(Bit#(64) _),
  function Action cache_0002_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0002(Bit#(64) _),
  function Action registerUL0002(Struct11 _),
  function ActionValue#(Bool) cache_0002_hasVictimSlot(),
  function Action makeEnq_parentChildren0002(Struct10 _),
  function ActionValue#(Bool) downLockable0002(Bit#(64) _),
  function ActionValue#(Bool) upLockable0002(Bit#(64) _),
  function ActionValue#(Struct31) cache_0002_readRs(),
  function ActionValue#(Struct2) deq_fifo000200(),
  function ActionValue#(Struct6) downLockRssFull0002(),
  function Action cache_0002_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00022()) (Module159);
    Reg#(Bit#(2)) rr0002 <- mkReg(unpack(0));
    Reg#(Struct30) prl0002 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0002 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0002 <- mkReg(unpack(0));
    Reg#(Struct5) wl0002 <- mkReg(unpack(0));

    rule rr_0002;let x_0 = (rr0002);
                 rr0002 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0002_1230;
        let x_0 = (prl0002);
        let x_1 = (crqrl0002);
        let x_2 = (crsrl0002);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00022();
        prl0002 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0002 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0002_readRq((x_3).addr);

    endrule

    rule rule_0002_1232;
        let x_0 = (prl0002);
        let x_1 = (crqrl0002);
        let x_2 = (crsrl0002);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0002();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0002 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0002 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0002_readRq((x_4).addr);

    endrule

    rule rule_0002_1231000200;
        let x_0 = (prl0002);
        let x_1 = (crqrl0002);
        let x_2 = (crsrl0002);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo000200();
        crqrl0002 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0002 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0002_readRq((x_3).addr);

    endrule

    rule rule_0002_456;
        let x_0 = (prl0002);
        let x_1 = (crqrl0002);
        let x_2 = (crsrl0002);
        let x_3 <- cache_0002_readRs();
        let x_4 = (rlc0002);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0002 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0002 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0002 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0002_00;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0002((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0002((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0002(x_17);
        let x_19 = (wl0002);
        when (! ((x_19).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0002_01;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0002((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0002_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0002(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0002(x_18);
        let x_20 = (wl0002);
        when (! ((x_20).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0002_020;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0002_writeRq(x_20);
        let x_22 <- releaseUL0002((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0002(x_23);
        let x_25 = (wl0002);
        when (! ((x_25).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_021;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0002_writeRq(x_20);
        let x_22 <- releaseUL0002((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0002(x_23);
        let x_25 = (wl0002);
        when (! ((x_25).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_03;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0002((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0002(x_19);
        let x_21 = (wl0002);
        when (! ((x_21).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_100;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0002((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0002((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0002_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0002(x_21);
        let x_23 = (wl0002);
        when (! ((x_23).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_101;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0002((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0002((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0002(x_19);
        let x_21 = (wl0002);
        when (! ((x_21).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_11;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0002((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0002_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0002(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0002(x_18);
        let x_20 = (wl0002);
        when (! ((x_20).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0002_12;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0002_writeRq(x_21);
        let x_23 <- releaseUL0002((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0002(x_24);
        let x_26 = (wl0002);
        when (! ((x_26).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_130;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0002((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0002(x_19);
        let x_21 = (wl0002);
        when (! ((x_21).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_131;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0002((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0002(x_19);
        let x_21 = (wl0002);
        when (! ((x_21).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0002_20;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        let x_4 <- cache_0002_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0002((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0002(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0002(x_16);
        let x_18 = (wl0002);
        when (! ((x_18).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0002_20, rule_0002_21" *)
    rule rule_0002_21;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        let x_4 <- cache_0002_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0002((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0002(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0002(x_16);
        let x_18 = (wl0002);
        when (! ((x_18).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0002_22;
        let x_0 = (rr0002);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0002);
        let x_2 = (crqrl0002);
        let x_3 = (crsrl0002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0002 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0002((x_11).addr);
        let x_18 = (wl0002);
        when (! ((x_18).wl_valid), noAction);
        wl0002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0002_removeVictim(x_19);
        let x_21 = (crqrl0002);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0002 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0002);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0002 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0002_7890;
        let x_0 = (wl0002);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0002 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0002_7891;
        let x_0 = (wl0002);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0002_writeRs();
        let x_2 = (prl0002);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0002 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0002);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0002 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0002);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0002 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0002 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module160;
endinterface


module mkModule160#(function ActionValue#(Struct31) cache_0003_writeRs(),
  function Action cache_0003_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0003_getVictim(),
  function Action releaseUL0003(Bit#(64) _),
  function Action cache_0003_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0003(Bit#(64) _),
  function Action registerUL0003(Struct11 _),
  function ActionValue#(Bool) cache_0003_hasVictimSlot(),
  function Action makeEnq_parentChildren0003(Struct10 _),
  function ActionValue#(Bool) downLockable0003(Bit#(64) _),
  function ActionValue#(Bool) upLockable0003(Bit#(64) _),
  function ActionValue#(Struct31) cache_0003_readRs(),
  function ActionValue#(Struct2) deq_fifo000300(),
  function ActionValue#(Struct6) downLockRssFull0003(),
  function Action cache_0003_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00032()) (Module160);
    Reg#(Bit#(2)) rr0003 <- mkReg(unpack(0));
    Reg#(Struct30) prl0003 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0003 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0003 <- mkReg(unpack(0));
    Reg#(Struct5) wl0003 <- mkReg(unpack(0));

    rule rr_0003;let x_0 = (rr0003);
                 rr0003 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0003_1230;
        let x_0 = (prl0003);
        let x_1 = (crqrl0003);
        let x_2 = (crsrl0003);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00032();
        prl0003 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0003 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0003_readRq((x_3).addr);

    endrule

    rule rule_0003_1232;
        let x_0 = (prl0003);
        let x_1 = (crqrl0003);
        let x_2 = (crsrl0003);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0003();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0003 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0003 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0003_readRq((x_4).addr);

    endrule

    rule rule_0003_1231000300;
        let x_0 = (prl0003);
        let x_1 = (crqrl0003);
        let x_2 = (crsrl0003);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo000300();
        crqrl0003 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0003 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0003_readRq((x_3).addr);

    endrule

    rule rule_0003_456;
        let x_0 = (prl0003);
        let x_1 = (crqrl0003);
        let x_2 = (crsrl0003);
        let x_3 <- cache_0003_readRs();
        let x_4 = (rlc0003);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0003 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0003 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0003 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0003_00;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0003((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0003((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0003(x_17);
        let x_19 = (wl0003);
        when (! ((x_19).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0003_01;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0003((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0003_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0003(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0003(x_18);
        let x_20 = (wl0003);
        when (! ((x_20).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0003_020;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0003_writeRq(x_20);
        let x_22 <- releaseUL0003((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0003(x_23);
        let x_25 = (wl0003);
        when (! ((x_25).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_021;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0003_writeRq(x_20);
        let x_22 <- releaseUL0003((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0003(x_23);
        let x_25 = (wl0003);
        when (! ((x_25).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_03;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0003((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0003(x_19);
        let x_21 = (wl0003);
        when (! ((x_21).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_100;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0003((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0003((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0003_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0003(x_21);
        let x_23 = (wl0003);
        when (! ((x_23).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_101;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0003((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0003((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0003(x_19);
        let x_21 = (wl0003);
        when (! ((x_21).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_11;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0003((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0003_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0003(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0003(x_18);
        let x_20 = (wl0003);
        when (! ((x_20).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0003_12;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0003_writeRq(x_21);
        let x_23 <- releaseUL0003((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0003(x_24);
        let x_26 = (wl0003);
        when (! ((x_26).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_130;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0003((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0003(x_19);
        let x_21 = (wl0003);
        when (! ((x_21).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_131;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0003((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0003(x_19);
        let x_21 = (wl0003);
        when (! ((x_21).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0003_20;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        let x_4 <- cache_0003_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0003((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0003(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0003(x_16);
        let x_18 = (wl0003);
        when (! ((x_18).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0003_20, rule_0003_21" *)
    rule rule_0003_21;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        let x_4 <- cache_0003_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0003((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0003(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0003(x_16);
        let x_18 = (wl0003);
        when (! ((x_18).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0003_22;
        let x_0 = (rr0003);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0003);
        let x_2 = (crqrl0003);
        let x_3 = (crsrl0003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0003 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0003((x_11).addr);
        let x_18 = (wl0003);
        when (! ((x_18).wl_valid), noAction);
        wl0003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0003_removeVictim(x_19);
        let x_21 = (crqrl0003);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0003 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0003);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0003 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0003_7890;
        let x_0 = (wl0003);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0003 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0003_7891;
        let x_0 = (wl0003);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0003_writeRs();
        let x_2 = (prl0003);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0003 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0003);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0003 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0003);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0003 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0003 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module161;
endinterface


module mkModule161#(function ActionValue#(Struct24) cache_001_writeRs(),
  function Action cache_001_removeVictim(Bit#(64) _),
  function ActionValue#(Struct24) cache_001_getVictim(),
  function Action transferUpDown001(Struct17 _),
  function Action releaseDL001(Bit#(64) _),
  function Action releaseUL001(Bit#(64) _),
  function ActionValue#(Struct15) upLockGet001(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00131(),
  function ActionValue#(Struct2) deq_fifo00121(),
  function ActionValue#(Struct2) deq_fifo00111(),
  function Action addRs001(Struct14 _),
  function ActionValue#(Struct6) downLockGet001(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00101(),
  function Action broadcast_parentChildren001(Struct13 _),
  function Action registerDL001(Struct12 _),
  function Action registerUL001(Struct11 _),
  function ActionValue#(Bool) cache_001_hasVictimSlot(),
  function Action makeEnq_parentChildren001(Struct10 _),
  function Action cache_001_writeRq(Struct24 _),
  function ActionValue#(Bool) downLockable001(Bit#(64) _),
  function ActionValue#(Bool) upLockable001(Bit#(64) _),
  function ActionValue#(Struct24) cache_001_readRs(),
  function ActionValue#(Struct2) deq_fifo00130(),
  function ActionValue#(Struct2) deq_fifo00120(),
  function ActionValue#(Struct2) deq_fifo00110(),
  function ActionValue#(Struct2) deq_fifo00100(),
  function ActionValue#(Struct6) downLockRssFull001(),
  function Action cache_001_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0012()) (Module161);
    Reg#(Bit#(2)) rr001 <- mkReg(unpack(0));
    Reg#(Struct23) prl001 <- mkReg(unpack(0));
    Reg#(Struct23) crqrl001 <- mkReg(unpack(0));
    Reg#(Struct23) crsrl001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc001 <- mkReg(unpack(0));
    Reg#(Struct5) wl001 <- mkReg(unpack(0));

    rule rr_001;let x_0 = (rr001);
                rr001 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_001_1230;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo0012();
        prl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc001 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_001_readRq((x_3).addr);

    endrule

    rule rule_001_1232;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull001();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc001 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_001_readRq((x_4).addr);

    endrule

    rule rule_001_123100100;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00100();
        crqrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc001 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_001_readRq((x_3).addr);

    endrule

    rule rule_001_123100110;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00110();
        crqrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h1), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc001 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_001_readRq((x_3).addr);

    endrule

    rule rule_001_123100120;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00120();
        crqrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h2), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc001 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_001_readRq((x_3).addr);

    endrule

    rule rule_001_123100130;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00130();
        crqrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h3), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc001 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_001_readRq((x_3).addr);

    endrule

    rule rule_001_456;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        let x_3 <- cache_001_readRs();
        let x_4 = (rlc001);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl001 <= Struct23 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl001 <= Struct23 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl001 <= Struct23 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_001_0000010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0010010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_010010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_030010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_100010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
        let x_23 = (wl001);
        when (! ((x_23).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_110010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_140010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_150010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        let x_17 <- broadcast_parentChildren001(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_250010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_26000010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_26010010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2610010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_270010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_280010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_2900010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2910010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2100010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2110010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_001_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 = (wl001);
        when (! ((x_24).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0400010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00101();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_0700010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00101();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16000010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00101();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16010010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00101();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110000010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00101();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110010010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00101();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110020010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00101();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_0000011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0010011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_010011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_030011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_100011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
        let x_23 = (wl001);
        when (! ((x_23).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_110011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_140011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_150011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        let x_17 <- broadcast_parentChildren001(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_250011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_26000011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_26010011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2610011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_270011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_280011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_2900011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2910011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2100011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2110011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_001_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 = (wl001);
        when (! ((x_24).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0400011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00111();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_0700011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00111();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16000011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00111();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16010011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00111();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110000011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00111();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110010011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00111();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110020011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00111();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_0000012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0010012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_010012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_030012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_100012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
        let x_23 = (wl001);
        when (! ((x_23).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_110012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_140012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_150012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        let x_17 <- broadcast_parentChildren001(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_250012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_26000012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_26010012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2610012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_270012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_280012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_2900012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2910012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2100012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2110012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_001_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 = (wl001);
        when (! ((x_24).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0400012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00121();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_0700012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00121();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16000012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00121();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16010012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00121();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110000012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00121();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110010012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00121();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110020012;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00121();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_0000013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0010013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_010013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_030013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_100013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren001(x_21);
        let x_23 = (wl001);
        when (! ((x_23).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_110013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_140013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_150013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((x_10).dir_sharers) &
        (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        let x_17 <- broadcast_parentChildren001(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_250013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_26000013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_26010013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2610013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_270013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_280013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_2900013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2910013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2100013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_001_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_21 <- makeEnq_parentChildren001(x_20);
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_2110013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_001_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 = (wl001);
        when (! ((x_24).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_0400013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00131();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_0700013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00131();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16000013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00131();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_16010013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00131();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110000013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00131();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110010013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00131();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_110020013;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        Struct24 x_4 =
        ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}));

        Bit#(64) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        let x_10 <- deq_fifo00131();
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_12 <- downLockGet001((x_10).addr);
        when ((x_12).valid, noAction);
        Struct7 x_13 = ((x_12).data);
        when (((x_10).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_13).dl_valid, noAction);
        when ((x_13).dl_rsb, noAction);
        when ((((x_13).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_10).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_14 = (x_10);
        let x_15 <- addRs001(Struct14 {r_dl_addr : (x_10).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_14});
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_020;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct24 x_22 = (Struct24 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_001_writeRq(x_22);
        let x_24 <- releaseUL001((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren001(x_25);
        let x_27 = (wl001);
        when (! ((x_27).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_021;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct24 x_22 = (Struct24 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_001_writeRq(x_22);
        let x_24 <- releaseUL001((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren001(x_25);
        let x_27 = (wl001);
        when (! ((x_27).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_041;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet001((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct24 x_18 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_st,
        mesi_dir_sharers : (((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_sharers) :
        (((Bit#(4))'(4'h1)) << ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_001_writeRq(x_21);
        let x_23 <- releaseDL001((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren001(x_24);
        let x_26 = (wl001);
        when (! ((x_26).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_05;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_10).dir_st))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_06;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_9))) && ((!
        (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_10).dir_st))))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h5)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_071;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet001((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct24 x_18 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0),
        dir_sharers : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (x_20).info_write, info : (x_20).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        let x_22 <- cache_001_writeRq(x_21);
        let x_23 <- releaseDL001((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren001(x_24);
        let x_26 = (wl001);
        when (! ((x_26).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_12;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((x_10).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))), noAction);

        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_001_writeRq(x_21);
        let x_23 <- releaseUL001((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren001(x_24);
        let x_26 = (wl001);
        when (! ((x_26).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_13;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))) ==
        ((Bit#(4))'(4'h0)))) && (((x_10).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = ((x_13).ul_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_18 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_19 <- cache_001_writeRq(x_18);
        let x_20 <- transferUpDown001(Struct17 {r_dl_addr : (x_11).addr,
        r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))});
        let x_21 <- broadcast_parentChildren001(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((x_17)[1:0]))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_16).addr, value : (Bit#(64))'(64'h0)}});
        let x_22 = (wl001);
        when (! ((x_22).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_161;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet001((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        let x_21 <- releaseDL001((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 = (wl001);
        when (! ((x_24).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_170;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_10).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_171;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_190;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h5)});
        let x_17 <- broadcast_parentChildren001(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_191;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h5)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_192;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL001(Struct12 {r_dl_rsb : (Bool)'(True),
        r_dl_msg : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h5)});
        let x_17 <- broadcast_parentChildren001(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value : (Bit#(64))'(64'h0)}});
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_11010;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet001((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        let x_21 <- releaseDL001((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 = (wl001);
        when (! ((x_24).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_11011;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct24 x_4 = ((x_3).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet001((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        let x_21 <- releaseDL001((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_23 <- makeEnq_parentChildren001(x_22);
        let x_24 = (wl001);
        when (! ((x_24).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_20;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        let x_4 <- cache_001_getVictim();
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_9))
        && ((x_9) < ((Bit#(3))'(3'h4)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        let x_15 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren001(x_16);
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_21;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        let x_4 <- cache_001_getVictim();
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when ((((x_10).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_8) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_9))) || (((x_8) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) && ((x_9) <
        ((Bit#(3))'(3'h3)))))), noAction);
        let x_15 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren001(x_16);
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_22;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL001((x_11).addr);
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_001_removeVictim(x_19);
        let x_21 = (crqrl001);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl001 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl001);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl001 <= Struct23 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    (* descending_urgency = "rule_001_23, rule_001_20, rule_001_21" *)
    rule rule_001_23;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        let x_4 <- cache_001_getVictim();
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((((x_9) == ((Bit#(3))'(3'h1))) && (! (((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_9) == ((Bit#(3))'(3'h2))) && ((x_8) ==
        ((Bool)'(False)))), noAction);
        let x_16 = (wl001);
        when (! ((x_16).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_17 = ((x_11).addr);
        let x_18 <- cache_001_removeVictim(x_17);
        let x_19 = (crqrl001);
        if ((((x_19).rl_valid) && ((x_19).rl_line_valid)) &&
        ((((x_19).rl_msg).addr) == (x_17))) begin

            crqrl001 <= Struct23 {rl_valid : (x_19).rl_valid, rl_cmidx :
            (x_19).rl_cmidx, rl_msg : (x_19).rl_msg, rl_line_valid :
            (x_19).rl_line_valid, rl_line : Struct24 {addr : x_17, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_21 = (crsrl001);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_17))) begin

            crsrl001 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_17, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 3'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_001_7890;
        let x_0 = (wl001);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl001 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_001_7891;
        let x_0 = (wl001);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_001_writeRs();
        let x_2 = (prl001);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl001);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl001);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl001 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module162;
endinterface


module mkModule162#(function ActionValue#(Struct31) cache_0010_writeRs(),
  function Action cache_0010_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0010_getVictim(),
  function Action releaseUL0010(Bit#(64) _),
  function Action cache_0010_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0010(Bit#(64) _),
  function Action registerUL0010(Struct11 _),
  function ActionValue#(Bool) cache_0010_hasVictimSlot(),
  function Action makeEnq_parentChildren0010(Struct10 _),
  function ActionValue#(Bool) downLockable0010(Bit#(64) _),
  function ActionValue#(Bool) upLockable0010(Bit#(64) _),
  function ActionValue#(Struct31) cache_0010_readRs(),
  function ActionValue#(Struct2) deq_fifo001000(),
  function ActionValue#(Struct6) downLockRssFull0010(),
  function Action cache_0010_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00102()) (Module162);
    Reg#(Bit#(2)) rr0010 <- mkReg(unpack(0));
    Reg#(Struct30) prl0010 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0010 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0010 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0010 <- mkReg(unpack(0));
    Reg#(Struct5) wl0010 <- mkReg(unpack(0));

    rule rr_0010;let x_0 = (rr0010);
                 rr0010 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0010_1230;
        let x_0 = (prl0010);
        let x_1 = (crqrl0010);
        let x_2 = (crsrl0010);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00102();
        prl0010 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0010 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0010_readRq((x_3).addr);

    endrule

    rule rule_0010_1232;
        let x_0 = (prl0010);
        let x_1 = (crqrl0010);
        let x_2 = (crsrl0010);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0010();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0010 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0010 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0010_readRq((x_4).addr);

    endrule

    rule rule_0010_1231001000;
        let x_0 = (prl0010);
        let x_1 = (crqrl0010);
        let x_2 = (crsrl0010);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo001000();
        crqrl0010 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0010 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0010_readRq((x_3).addr);

    endrule

    rule rule_0010_456;
        let x_0 = (prl0010);
        let x_1 = (crqrl0010);
        let x_2 = (crsrl0010);
        let x_3 <- cache_0010_readRs();
        let x_4 = (rlc0010);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0010 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0010 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0010 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0010_00;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0010((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0010((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0010(x_17);
        let x_19 = (wl0010);
        when (! ((x_19).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0010_01;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0010((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0010_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0010(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0010(x_18);
        let x_20 = (wl0010);
        when (! ((x_20).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0010_020;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0010((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0010((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0010_writeRq(x_20);
        let x_22 <- releaseUL0010((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0010(x_23);
        let x_25 = (wl0010);
        when (! ((x_25).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_021;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0010((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0010((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0010_writeRq(x_20);
        let x_22 <- releaseUL0010((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0010(x_23);
        let x_25 = (wl0010);
        when (! ((x_25).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_03;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0010((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0010_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0010(x_19);
        let x_21 = (wl0010);
        when (! ((x_21).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_100;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0010((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0010((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0010_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0010(x_21);
        let x_23 = (wl0010);
        when (! ((x_23).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_101;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0010((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0010((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0010_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0010(x_19);
        let x_21 = (wl0010);
        when (! ((x_21).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_11;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0010((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0010_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0010(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0010(x_18);
        let x_20 = (wl0010);
        when (! ((x_20).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0010_12;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0010((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0010((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0010_writeRq(x_21);
        let x_23 <- releaseUL0010((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0010(x_24);
        let x_26 = (wl0010);
        when (! ((x_26).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_130;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0010((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0010_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0010(x_19);
        let x_21 = (wl0010);
        when (! ((x_21).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_131;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0010((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0010_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0010(x_19);
        let x_21 = (wl0010);
        when (! ((x_21).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0010_20;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        let x_4 <- cache_0010_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0010((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0010(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0010(x_16);
        let x_18 = (wl0010);
        when (! ((x_18).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0010_20, rule_0010_21" *)
    rule rule_0010_21;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        let x_4 <- cache_0010_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0010((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0010(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0010(x_16);
        let x_18 = (wl0010);
        when (! ((x_18).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0010_22;
        let x_0 = (rr0010);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0010);
        let x_2 = (crqrl0010);
        let x_3 = (crsrl0010);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0010((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0010((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0010 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0010((x_11).addr);
        let x_18 = (wl0010);
        when (! ((x_18).wl_valid), noAction);
        wl0010 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0010_removeVictim(x_19);
        let x_21 = (crqrl0010);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0010 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0010);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0010 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0010_7890;
        let x_0 = (wl0010);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0010 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0010_7891;
        let x_0 = (wl0010);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0010_writeRs();
        let x_2 = (prl0010);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0010 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0010);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0010 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0010);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0010 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0010 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module163;
endinterface


module mkModule163#(function ActionValue#(Struct31) cache_0011_writeRs(),
  function Action cache_0011_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0011_getVictim(),
  function Action releaseUL0011(Bit#(64) _),
  function Action cache_0011_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0011(Bit#(64) _),
  function Action registerUL0011(Struct11 _),
  function ActionValue#(Bool) cache_0011_hasVictimSlot(),
  function Action makeEnq_parentChildren0011(Struct10 _),
  function ActionValue#(Bool) downLockable0011(Bit#(64) _),
  function ActionValue#(Bool) upLockable0011(Bit#(64) _),
  function ActionValue#(Struct31) cache_0011_readRs(),
  function ActionValue#(Struct2) deq_fifo001100(),
  function ActionValue#(Struct6) downLockRssFull0011(),
  function Action cache_0011_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00112()) (Module163);
    Reg#(Bit#(2)) rr0011 <- mkReg(unpack(0));
    Reg#(Struct30) prl0011 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0011 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0011 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0011 <- mkReg(unpack(0));
    Reg#(Struct5) wl0011 <- mkReg(unpack(0));

    rule rr_0011;let x_0 = (rr0011);
                 rr0011 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0011_1230;
        let x_0 = (prl0011);
        let x_1 = (crqrl0011);
        let x_2 = (crsrl0011);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00112();
        prl0011 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0011 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0011_readRq((x_3).addr);

    endrule

    rule rule_0011_1232;
        let x_0 = (prl0011);
        let x_1 = (crqrl0011);
        let x_2 = (crsrl0011);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0011();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0011 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0011 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0011_readRq((x_4).addr);

    endrule

    rule rule_0011_1231001100;
        let x_0 = (prl0011);
        let x_1 = (crqrl0011);
        let x_2 = (crsrl0011);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo001100();
        crqrl0011 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0011 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0011_readRq((x_3).addr);

    endrule

    rule rule_0011_456;
        let x_0 = (prl0011);
        let x_1 = (crqrl0011);
        let x_2 = (crsrl0011);
        let x_3 <- cache_0011_readRs();
        let x_4 = (rlc0011);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0011 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0011 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0011 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0011_00;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0011((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0011((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0011(x_17);
        let x_19 = (wl0011);
        when (! ((x_19).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0011_01;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0011((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0011_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0011(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0011(x_18);
        let x_20 = (wl0011);
        when (! ((x_20).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0011_020;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0011((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0011((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0011_writeRq(x_20);
        let x_22 <- releaseUL0011((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0011(x_23);
        let x_25 = (wl0011);
        when (! ((x_25).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_021;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0011((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0011((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0011_writeRq(x_20);
        let x_22 <- releaseUL0011((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0011(x_23);
        let x_25 = (wl0011);
        when (! ((x_25).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_03;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0011((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0011_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0011(x_19);
        let x_21 = (wl0011);
        when (! ((x_21).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_100;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0011((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0011((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0011_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0011(x_21);
        let x_23 = (wl0011);
        when (! ((x_23).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_101;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0011((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0011((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0011_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0011(x_19);
        let x_21 = (wl0011);
        when (! ((x_21).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_11;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0011((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0011_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0011(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0011(x_18);
        let x_20 = (wl0011);
        when (! ((x_20).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0011_12;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0011((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0011((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0011_writeRq(x_21);
        let x_23 <- releaseUL0011((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0011(x_24);
        let x_26 = (wl0011);
        when (! ((x_26).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_130;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0011((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0011_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0011(x_19);
        let x_21 = (wl0011);
        when (! ((x_21).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_131;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0011((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0011_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0011(x_19);
        let x_21 = (wl0011);
        when (! ((x_21).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0011_20;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        let x_4 <- cache_0011_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0011((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0011(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0011(x_16);
        let x_18 = (wl0011);
        when (! ((x_18).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0011_20, rule_0011_21" *)
    rule rule_0011_21;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        let x_4 <- cache_0011_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0011((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0011(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0011(x_16);
        let x_18 = (wl0011);
        when (! ((x_18).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0011_22;
        let x_0 = (rr0011);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0011);
        let x_2 = (crqrl0011);
        let x_3 = (crsrl0011);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0011((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0011((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0011 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0011((x_11).addr);
        let x_18 = (wl0011);
        when (! ((x_18).wl_valid), noAction);
        wl0011 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0011_removeVictim(x_19);
        let x_21 = (crqrl0011);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0011 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0011);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0011 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0011_7890;
        let x_0 = (wl0011);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0011 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0011_7891;
        let x_0 = (wl0011);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0011_writeRs();
        let x_2 = (prl0011);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0011 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0011);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0011 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0011);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0011 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0011 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module164;
endinterface


module mkModule164#(function ActionValue#(Struct31) cache_0012_writeRs(),
  function Action cache_0012_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0012_getVictim(),
  function Action releaseUL0012(Bit#(64) _),
  function Action cache_0012_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0012(Bit#(64) _),
  function Action registerUL0012(Struct11 _),
  function ActionValue#(Bool) cache_0012_hasVictimSlot(),
  function Action makeEnq_parentChildren0012(Struct10 _),
  function ActionValue#(Bool) downLockable0012(Bit#(64) _),
  function ActionValue#(Bool) upLockable0012(Bit#(64) _),
  function ActionValue#(Struct31) cache_0012_readRs(),
  function ActionValue#(Struct2) deq_fifo001200(),
  function ActionValue#(Struct6) downLockRssFull0012(),
  function Action cache_0012_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00122()) (Module164);
    Reg#(Bit#(2)) rr0012 <- mkReg(unpack(0));
    Reg#(Struct30) prl0012 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0012 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0012 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0012 <- mkReg(unpack(0));
    Reg#(Struct5) wl0012 <- mkReg(unpack(0));

    rule rr_0012;let x_0 = (rr0012);
                 rr0012 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0012_1230;
        let x_0 = (prl0012);
        let x_1 = (crqrl0012);
        let x_2 = (crsrl0012);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00122();
        prl0012 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0012 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0012_readRq((x_3).addr);

    endrule

    rule rule_0012_1232;
        let x_0 = (prl0012);
        let x_1 = (crqrl0012);
        let x_2 = (crsrl0012);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0012();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0012 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0012 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0012_readRq((x_4).addr);

    endrule

    rule rule_0012_1231001200;
        let x_0 = (prl0012);
        let x_1 = (crqrl0012);
        let x_2 = (crsrl0012);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo001200();
        crqrl0012 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0012 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0012_readRq((x_3).addr);

    endrule

    rule rule_0012_456;
        let x_0 = (prl0012);
        let x_1 = (crqrl0012);
        let x_2 = (crsrl0012);
        let x_3 <- cache_0012_readRs();
        let x_4 = (rlc0012);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0012 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0012 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0012 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0012_00;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0012((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0012((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0012(x_17);
        let x_19 = (wl0012);
        when (! ((x_19).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0012_01;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0012((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0012_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0012(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0012(x_18);
        let x_20 = (wl0012);
        when (! ((x_20).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0012_020;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0012((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0012((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0012_writeRq(x_20);
        let x_22 <- releaseUL0012((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0012(x_23);
        let x_25 = (wl0012);
        when (! ((x_25).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_021;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0012((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0012((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0012_writeRq(x_20);
        let x_22 <- releaseUL0012((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0012(x_23);
        let x_25 = (wl0012);
        when (! ((x_25).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_03;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0012((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0012_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0012(x_19);
        let x_21 = (wl0012);
        when (! ((x_21).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_100;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0012((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0012((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0012_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0012(x_21);
        let x_23 = (wl0012);
        when (! ((x_23).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_101;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0012((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0012((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0012_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0012(x_19);
        let x_21 = (wl0012);
        when (! ((x_21).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_11;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0012((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0012_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0012(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0012(x_18);
        let x_20 = (wl0012);
        when (! ((x_20).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0012_12;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0012((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0012((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0012_writeRq(x_21);
        let x_23 <- releaseUL0012((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0012(x_24);
        let x_26 = (wl0012);
        when (! ((x_26).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_130;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0012((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0012_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0012(x_19);
        let x_21 = (wl0012);
        when (! ((x_21).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_131;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0012((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0012_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0012(x_19);
        let x_21 = (wl0012);
        when (! ((x_21).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0012_20;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        let x_4 <- cache_0012_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0012((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0012(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0012(x_16);
        let x_18 = (wl0012);
        when (! ((x_18).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0012_20, rule_0012_21" *)
    rule rule_0012_21;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        let x_4 <- cache_0012_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0012((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0012(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0012(x_16);
        let x_18 = (wl0012);
        when (! ((x_18).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0012_22;
        let x_0 = (rr0012);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0012);
        let x_2 = (crqrl0012);
        let x_3 = (crsrl0012);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0012((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0012((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0012 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0012((x_11).addr);
        let x_18 = (wl0012);
        when (! ((x_18).wl_valid), noAction);
        wl0012 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0012_removeVictim(x_19);
        let x_21 = (crqrl0012);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0012 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0012);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0012 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0012_7890;
        let x_0 = (wl0012);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0012 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0012_7891;
        let x_0 = (wl0012);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0012_writeRs();
        let x_2 = (prl0012);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0012 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0012);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0012 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0012);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0012 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0012 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module165;
endinterface


module mkModule165#(function ActionValue#(Struct31) cache_0013_writeRs(),
  function Action cache_0013_removeVictim(Bit#(64) _),
  function ActionValue#(Struct31) cache_0013_getVictim(),
  function Action releaseUL0013(Bit#(64) _),
  function Action cache_0013_writeRq(Struct31 _),
  function ActionValue#(Struct15) upLockGet0013(Bit#(64) _),
  function Action registerUL0013(Struct11 _),
  function ActionValue#(Bool) cache_0013_hasVictimSlot(),
  function Action makeEnq_parentChildren0013(Struct10 _),
  function ActionValue#(Bool) downLockable0013(Bit#(64) _),
  function ActionValue#(Bool) upLockable0013(Bit#(64) _),
  function ActionValue#(Struct31) cache_0013_readRs(),
  function ActionValue#(Struct2) deq_fifo001300(),
  function ActionValue#(Struct6) downLockRssFull0013(),
  function Action cache_0013_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo00132()) (Module165);
    Reg#(Bit#(2)) rr0013 <- mkReg(unpack(0));
    Reg#(Struct30) prl0013 <- mkReg(unpack(0));
    Reg#(Struct30) crqrl0013 <- mkReg(unpack(0));
    Reg#(Struct30) crsrl0013 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc0013 <- mkReg(unpack(0));
    Reg#(Struct5) wl0013 <- mkReg(unpack(0));

    rule rr_0013;let x_0 = (rr0013);
                 rr0013 <= (x_0) + ((Bit#(2))'(2'h1));

    endrule

    rule rule_0013_1230;
        let x_0 = (prl0013);
        let x_1 = (crqrl0013);
        let x_2 = (crsrl0013);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo00132();
        prl0013 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0013 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_0013_readRq((x_3).addr);

    endrule

    rule rule_0013_1232;
        let x_0 = (prl0013);
        let x_1 = (crqrl0013);
        let x_2 = (crsrl0013);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull0013();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl0013 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0013 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_0013_readRq((x_4).addr);

    endrule

    rule rule_0013_1231001300;
        let x_0 = (prl0013);
        let x_1 = (crqrl0013);
        let x_2 = (crsrl0013);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo001300();
        crqrl0013 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})};

        rlc0013 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_0013_readRq((x_3).addr);

    endrule

    rule rule_0013_456;
        let x_0 = (prl0013);
        let x_1 = (crqrl0013);
        let x_2 = (crsrl0013);
        let x_3 <- cache_0013_readRs();
        let x_4 = (rlc0013);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl0013 <= Struct30 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl0013 <= Struct30 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl0013 <= Struct30 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_0013_00;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0013((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0013((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren0013(x_17);
        let x_19 = (wl0013);
        when (! ((x_19).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0013_01;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0013((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0013_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0013(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0013(x_18);
        let x_20 = (wl0013);
        when (! ((x_20).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0013_020;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0013((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0013((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0013_writeRq(x_20);
        let x_22 <- releaseUL0013((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0013(x_23);
        let x_25 = (wl0013);
        when (! ((x_25).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_021;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0013((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0013((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_0013_writeRq(x_20);
        let x_22 <- releaseUL0013((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren0013(x_23);
        let x_25 = (wl0013);
        when (! ((x_25).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_03;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0013((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0013_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren0013(x_19);
        let x_21 = (wl0013);
        when (! ((x_21).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_100;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0013((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0013((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct31 x_18 = (Struct31 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct31 x_19 = (Struct31 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_0013_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_22 <- makeEnq_parentChildren0013(x_21);
        let x_23 = (wl0013);
        when (! ((x_23).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_101;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0013((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable0013((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct31 x_17 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_0013_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0013(x_19);
        let x_21 = (wl0013);
        when (! ((x_21).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_11;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct31 x_4 = ((x_2).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0013((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_0013_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL0013(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_19 <- makeEnq_parentChildren0013(x_18);
        let x_20 = (wl0013);
        when (! ((x_20).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0013_12;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0013((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0013((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct31 x_19 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct31 x_20 = (Struct31 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct31 x_21 = (Struct31 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_0013_writeRq(x_21);
        let x_23 <- releaseUL0013((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_25 <- makeEnq_parentChildren0013(x_24);
        let x_26 = (wl0013);
        when (! ((x_26).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_130;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0013((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0013_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0013(x_19);
        let x_21 = (wl0013);
        when (! ((x_21).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_131;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable0013((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_15 = (x_11);
        Struct31 x_16 = (Struct31 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct31 x_17 = (Struct31 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_0013_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Bit#(64))'(64'h0)}});
        let x_20 <- makeEnq_parentChildren0013(x_19);
        let x_21 = (wl0013);
        when (! ((x_21).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_0013_20;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        let x_4 <- cache_0013_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0013((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_9)) &&
        ((x_9) < ((Bit#(3))'(3'h4)))), noAction);
        let x_15 <- registerUL0013(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_11).addr, value
        : (Bit#(64))'(64'h0)}});
        let x_17 <- makeEnq_parentChildren0013(x_16);
        let x_18 = (wl0013);
        when (! ((x_18).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_0013_20, rule_0013_21" *)
    rule rule_0013_21;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h3)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        let x_4 <- cache_0013_getVictim();
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_5).addr, value : (Bit#(64))'(64'h0)});

        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable0013((x_11).addr);
        when (x_14, noAction);
        when (((Bit#(3))'(3'h0)) < (x_9), noAction);
        let x_15 <- registerUL0013(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_11, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_16 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_11).addr, value
        : x_6}});
        let x_17 <- makeEnq_parentChildren0013(x_16);
        let x_18 = (wl0013);
        when (! ((x_18).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_0013_22;
        let x_0 = (rr0013);
        when ((x_0) == ((Bit#(2))'(2'h0)), noAction);
        let x_1 = (prl0013);
        let x_2 = (crqrl0013);
        let x_3 = (crsrl0013);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct31 x_4 = ((x_1).rl_line);
        Struct31 x_5 = (Struct31 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Bit#(64) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet0013((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable0013((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl0013 <=
        (Struct30)'(Struct30 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: 64'h0}, rl_line_valid: False, rl_line: Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL0013((x_11).addr);
        let x_18 = (wl0013);
        when (! ((x_18).wl_valid), noAction);
        wl0013 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_0013_removeVictim(x_19);
        let x_21 = (crqrl0013);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl0013 <= Struct30 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end
        let x_23 = (crsrl0013);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl0013 <= Struct30 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct31 {addr : x_19, info_hit :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_hit,
            info_way :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_way,
            info_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info_write,
            info :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).info,
            value_write :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value_write,
            value :
            ((Struct31)'(Struct31 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: 64'h0})).value}};


        end else begin

        end

    endrule

    rule rule_0013_7890;
        let x_0 = (wl0013);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl0013 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_0013_7891;
        let x_0 = (wl0013);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_0013_writeRs();
        let x_2 = (prl0013);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl0013 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl0013);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl0013 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl0013);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl0013 <= Struct30 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl0013 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule


interface CC;
    method Action mem_enq_rq_0 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_0 ();
    method Action mem_enq_rq_1 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_1 ();
    method Action mem_enq_rq_2 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_2 ();
    method Action mem_enq_rq_3 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_3 ();
    method Action mem_enq_rq_4 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_4 ();
    method Action mem_enq_rq_5 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_5 ();
    method Action mem_enq_rq_6 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_6 ();
    method Action mem_enq_rq_7 (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs_7 ();

    method Bool isInit ();
endinterface

module mkCC#(function ActionValue#(Struct2) deq_fifo002(),
  function Action enq_fifo0022(Struct2 _),
  function Action enq_fifo0032(Struct2 _),
  function Action enq_fifo001(Struct2 _),
  function Action enq_fifo000(Struct2 _)) (CC);
    Module1 m1 <- mkModule1 ();
    Module2 m2 <- mkModule2 ();
    Module3 m3 <- mkModule3 ();
    Module4 m4 <- mkModule4 ();
    Module5 m5 <- mkModule5 ();
    Module6 m6 <- mkModule6 ();
    Module7 m7 <- mkModule7 ();
    Module8 m8 <- mkModule8 ();
    Module9 m9 <- mkModule9 ();
    Module10 m10 <- mkModule10 ();
    Module11 m11 <- mkModule11 ();
    Module12 m12 <- mkModule12 ();
    Module13 m13 <- mkModule13 ();
    Module14 m14 <- mkModule14 ();
    Module15 m15 <- mkModule15 ();
    Module16 m16 <- mkModule16 ();
    Module17 m17 <- mkModule17 ();
    Module18 m18 <- mkModule18 ();
    Module19 m19 <- mkModule19 ();
    Module20 m20 <- mkModule20 ();
    Module21 m21 <- mkModule21 ();
    Module22 m22 <- mkModule22 ();
    Module23 m23 <- mkModule23 ();
    Module24 m24 <- mkModule24 ();
    Module25 m25 <- mkModule25 ();
    Module26 m26 <- mkModule26 ();
    Module27 m27 <- mkModule27 ();
    Module28 m28 <- mkModule28 ();
    Module29 m29 <- mkModule29 ();
    Module30 m30 <- mkModule30 ();
    Module31 m31 <- mkModule31 ();
    Module32 m32 <- mkModule32 ();
    Module33 m33 <- mkModule33 ();
    Module34 m34 <- mkModule34 ();
    Module35 m35 <- mkModule35 ();
    Module36 m36 <- mkModule36 ();
    Module37 m37 <- mkModule37 ();
    Module38 m38 <- mkModule38 ();
    Module39 m39 <- mkModule39 ();
    Module40 m40 <- mkModule40 ();
    Module41 m41 <- mkModule41 ();
    Module42 m42 <- mkModule42 ();
    Module43 m43 <- mkModule43 ();
    Module44 m44 <- mkModule44 ();
    Module45 m45 <- mkModule45 ();
    Module46 m46 <- mkModule46 ();
    Module47 m47 <- mkModule47 ();
    Module48 m48 <- mkModule48 ();
    Module49 m49 <- mkModule49 ();
    Module50 m50 <- mkModule50 ();
    Module51 m51 <- mkModule51 ();
    Module52 m52 <- mkModule52 ();
    Module53 m53 <- mkModule53 ();
    Module54 m54 <- mkModule54 ();
    Module55 m55 <- mkModule55 ();
    Module56 m56 <- mkModule56 ();
    Module57 m57 <- mkModule57 ();
    Module58 m58 <- mkModule58 ();
    Module59 m59 <- mkModule59 ();
    Module60 m60 <- mkModule60 ();
    Module61 m61 <- mkModule61 ();
    Module62 m62 <- mkModule62 ();
    Module63 m63 <- mkModule63 ();
    Module64 m64 <- mkModule64 ();
    Module65 m65 <- mkModule65 ();
    Module66 m66 <- mkModule66 ();
    Module67 m67 <- mkModule67 ();
    Module68 m68 <- mkModule68 ();
    Module69 m69 <- mkModule69 ();
    Module70 m70 <- mkModule70 ();
    Module71 m71 <- mkModule71 ();
    Module72 m72 <- mkModule72 ();
    Module73 m73 <- mkModule73 ();
    Module74 m74 <- mkModule74 ();
    Module75 m75 <- mkModule75 ();
    Module76 m76 <- mkModule76 ();
    Module77 m77 <- mkModule77 ();
    Module78 m78 <- mkModule78 ();
    Module79 m79 <- mkModule79 ();
    Module80 m80 <- mkModule80 ();
    Module81 m81 <- mkModule81 ();
    Module82 m82 <- mkModule82 ();
    Module83 m83 <- mkModule83 ();
    Module84 m84 <- mkModule84 ();
    Module85 m85 <- mkModule85 ();
    Module86 m86 <- mkModule86 ();
    Module87 m87 <- mkModule87 ();
    Module88 m88 <- mkModule88 ();
    Module89 m89 <- mkModule89 ();
    Module90 m90 <- mkModule90 ();
    Module91 m91 <- mkModule91 ();
    Module92 m92 <- mkModule92 ();
    Module93 m93 <- mkModule93 ();
    Module94 m94 <- mkModule94 ();
    Module95 m95 <- mkModule95 ();
    Module96 m96 <- mkModule96 ();
    Module97 m97 <- mkModule97 ();
    Module98 m98 <- mkModule98 ();
    Module99 m99 <- mkModule99 ();
    Module100 m100 <- mkModule100 ();
    Module101 m101 <- mkModule101 ();
    Module102 m102 <- mkModule102 ();
    Module103 m103 <- mkModule103 ();
    Module104 m104 <- mkModule104 ();
    Module105 m105 <- mkModule105 ();
    Module106 m106 <- mkModule106 ();
    Module107 m107 <- mkModule107 ();
    Module108 m108 <- mkModule108 ();
    Module109 m109 <- mkModule109 ();
    Module110 m110 <- mkModule110 ();
    Module111 m111 <- mkModule111 ();
    Module112 m112 <- mkModule112 ();
    Module113 m113 <- mkModule113 ();
    Module114 m114 <- mkModule114 ();
    Module115 m115 <- mkModule115 ();
    Module116 m116 <- mkModule116 ();
    Module117 m117 <- mkModule117 ();
    Module118 m118 <- mkModule118 ();
    Module119 m119 <- mkModule119 ();
    Module120 m120 <- mkModule120 ();
    Module121 m121 <- mkModule121 ();
    Module122 m122 <- mkModule122 ();
    Module123 m123 <- mkModule123 ();
    Module124 m124 <- mkModule124 ();
    Module125 m125 <- mkModule125 ();
    Module126 m126 <- mkModule126 ();
    Module127 m127 <- mkModule127 ();
    Module128 m128 <- mkModule128 ();
    Module129 m129 <- mkModule129 ();
    Module130 m130 <- mkModule130 ();
    Module131 m131 <- mkModule131 ();
    Module132 m132 <- mkModule132 ();
    Module133 m133 <- mkModule133 (m1.putRq_infoRam_00_15,
    m2.putRq_infoRam_00_14, m3.putRq_infoRam_00_13, m4.putRq_infoRam_00_12,
    m5.putRq_infoRam_00_11, m6.putRq_infoRam_00_10, m7.putRq_infoRam_00_9,
    m8.putRq_infoRam_00_8, m9.putRq_infoRam_00_7, m10.putRq_infoRam_00_6,
    m11.putRq_infoRam_00_5, m12.putRq_infoRam_00_4, m13.putRq_infoRam_00_3,
    m14.putRq_infoRam_00_2, m15.putRq_infoRam_00_1, m16.putRq_infoRam_00_0,
    m17.getRs_dataRam_00, m17.putRq_dataRam_00, m1.getRs_infoRam_00_15,
    m2.getRs_infoRam_00_14, m3.getRs_infoRam_00_13, m4.getRs_infoRam_00_12,
    m5.getRs_infoRam_00_11, m6.getRs_infoRam_00_10, m7.getRs_infoRam_00_9,
    m8.getRs_infoRam_00_8, m9.getRs_infoRam_00_7, m10.getRs_infoRam_00_6,
    m11.getRs_infoRam_00_5, m12.getRs_infoRam_00_4, m13.getRs_infoRam_00_3,
    m14.getRs_infoRam_00_2, m15.getRs_infoRam_00_1, m16.getRs_infoRam_00_0);

    Module134 m134 <- mkModule134 (m31.enq_fifo0002, m88.enq_fifo0012,
    enq_fifo0022, enq_fifo0032, enq_fifo001, enq_fifo000);
    Module135 m135 <- mkModule135 (m19.putRq_infoRam_000_7,
    m20.putRq_infoRam_000_6, m21.putRq_infoRam_000_5,
    m22.putRq_infoRam_000_4, m23.putRq_infoRam_000_3,
    m24.putRq_infoRam_000_2, m25.putRq_infoRam_000_1,
    m26.putRq_infoRam_000_0, m27.getRs_dataRam_000, m27.putRq_dataRam_000,
    m19.getRs_infoRam_000_7, m20.getRs_infoRam_000_6,
    m21.getRs_infoRam_000_5, m22.getRs_infoRam_000_4,
    m23.getRs_infoRam_000_3, m24.getRs_infoRam_000_2,
    m25.getRs_infoRam_000_1, m26.getRs_infoRam_000_0);
    Module136 m136 <- mkModule136 (m40.enq_fifo00002, m51.enq_fifo00012,
    m62.enq_fifo00022, m73.enq_fifo00032, m30.enq_fifo0001,
    m29.enq_fifo0000);
    Module137 m137 <- mkModule137 (m32.putRq_infoRam_0000_3,
    m33.putRq_infoRam_0000_2, m34.putRq_infoRam_0000_1,
    m35.putRq_infoRam_0000_0, m36.getRs_dataRam_0000, m36.putRq_dataRam_0000,
    m32.getRs_infoRam_0000_3, m33.getRs_infoRam_0000_2,
    m34.getRs_infoRam_0000_1, m35.getRs_infoRam_0000_0);
    Module138 m138 <- mkModule138 (m42.enq_fifo000002, m39.enq_fifo00001,
    m38.enq_fifo00000);
    Module139 m139 <- mkModule139 (m43.putRq_infoRam_0001_3,
    m44.putRq_infoRam_0001_2, m45.putRq_infoRam_0001_1,
    m46.putRq_infoRam_0001_0, m47.getRs_dataRam_0001, m47.putRq_dataRam_0001,
    m43.getRs_infoRam_0001_3, m44.getRs_infoRam_0001_2,
    m45.getRs_infoRam_0001_1, m46.getRs_infoRam_0001_0);
    Module140 m140 <- mkModule140 (m53.enq_fifo000102, m50.enq_fifo00011,
    m49.enq_fifo00010);
    Module141 m141 <- mkModule141 (m54.putRq_infoRam_0002_3,
    m55.putRq_infoRam_0002_2, m56.putRq_infoRam_0002_1,
    m57.putRq_infoRam_0002_0, m58.getRs_dataRam_0002, m58.putRq_dataRam_0002,
    m54.getRs_infoRam_0002_3, m55.getRs_infoRam_0002_2,
    m56.getRs_infoRam_0002_1, m57.getRs_infoRam_0002_0);
    Module142 m142 <- mkModule142 (m64.enq_fifo000202, m61.enq_fifo00021,
    m60.enq_fifo00020);
    Module143 m143 <- mkModule143 (m65.putRq_infoRam_0003_3,
    m66.putRq_infoRam_0003_2, m67.putRq_infoRam_0003_1,
    m68.putRq_infoRam_0003_0, m69.getRs_dataRam_0003, m69.putRq_dataRam_0003,
    m65.getRs_infoRam_0003_3, m66.getRs_infoRam_0003_2,
    m67.getRs_infoRam_0003_1, m68.getRs_infoRam_0003_0);
    Module144 m144 <- mkModule144 (m75.enq_fifo000302, m72.enq_fifo00031,
    m71.enq_fifo00030);
    Module145 m145 <- mkModule145 (m76.putRq_infoRam_001_7,
    m77.putRq_infoRam_001_6, m78.putRq_infoRam_001_5,
    m79.putRq_infoRam_001_4, m80.putRq_infoRam_001_3,
    m81.putRq_infoRam_001_2, m82.putRq_infoRam_001_1,
    m83.putRq_infoRam_001_0, m84.getRs_dataRam_001, m84.putRq_dataRam_001,
    m76.getRs_infoRam_001_7, m77.getRs_infoRam_001_6,
    m78.getRs_infoRam_001_5, m79.getRs_infoRam_001_4,
    m80.getRs_infoRam_001_3, m81.getRs_infoRam_001_2,
    m82.getRs_infoRam_001_1, m83.getRs_infoRam_001_0);
    Module146 m146 <- mkModule146 (m97.enq_fifo00102, m108.enq_fifo00112,
    m119.enq_fifo00122, m130.enq_fifo00132, m87.enq_fifo0011,
    m86.enq_fifo0010);
    Module147 m147 <- mkModule147 (m89.putRq_infoRam_0010_3,
    m90.putRq_infoRam_0010_2, m91.putRq_infoRam_0010_1,
    m92.putRq_infoRam_0010_0, m93.getRs_dataRam_0010, m93.putRq_dataRam_0010,
    m89.getRs_infoRam_0010_3, m90.getRs_infoRam_0010_2,
    m91.getRs_infoRam_0010_1, m92.getRs_infoRam_0010_0);
    Module148 m148 <- mkModule148 (m99.enq_fifo001002, m96.enq_fifo00101,
    m95.enq_fifo00100);
    Module149 m149 <- mkModule149 (m100.putRq_infoRam_0011_3,
    m101.putRq_infoRam_0011_2, m102.putRq_infoRam_0011_1,
    m103.putRq_infoRam_0011_0, m104.getRs_dataRam_0011,
    m104.putRq_dataRam_0011, m100.getRs_infoRam_0011_3,
    m101.getRs_infoRam_0011_2, m102.getRs_infoRam_0011_1,
    m103.getRs_infoRam_0011_0);
    Module150 m150 <- mkModule150 (m110.enq_fifo001102, m107.enq_fifo00111,
    m106.enq_fifo00110);
    Module151 m151 <- mkModule151 (m111.putRq_infoRam_0012_3,
    m112.putRq_infoRam_0012_2, m113.putRq_infoRam_0012_1,
    m114.putRq_infoRam_0012_0, m115.getRs_dataRam_0012,
    m115.putRq_dataRam_0012, m111.getRs_infoRam_0012_3,
    m112.getRs_infoRam_0012_2, m113.getRs_infoRam_0012_1,
    m114.getRs_infoRam_0012_0);
    Module152 m152 <- mkModule152 (m121.enq_fifo001202, m118.enq_fifo00121,
    m117.enq_fifo00120);
    Module153 m153 <- mkModule153 (m122.putRq_infoRam_0013_3,
    m123.putRq_infoRam_0013_2, m124.putRq_infoRam_0013_1,
    m125.putRq_infoRam_0013_0, m126.getRs_dataRam_0013,
    m126.putRq_dataRam_0013, m122.getRs_infoRam_0013_3,
    m123.getRs_infoRam_0013_2, m124.getRs_infoRam_0013_1,
    m125.getRs_infoRam_0013_0);
    Module154 m154 <- mkModule154 (m132.enq_fifo001302, m129.enq_fifo00131,
    m128.enq_fifo00130);
    Module155 m155 <- mkModule155 (m133.cache_00_writeRs,
    m133.cache_00_removeVictim, m133.cache_00_getVictim,
    m18.transferUpDown00, m18.releaseDL00, m18.releaseUL00, m18.upLockGet00,
    m87.deq_fifo0011, m18.addRs00, m18.downLockGet00, m30.deq_fifo0001,
    m134.broadcast_parentChildren00, m18.registerDL00, m18.registerUL00,
    m133.cache_00_hasVictimSlot, m134.makeEnq_parentChildren00,
    m133.cache_00_writeRq, m18.downLockable00, m18.upLockable00,
    m133.cache_00_readRs, m86.deq_fifo0010, m29.deq_fifo0000,
    m18.downLockRssFull00, m133.cache_00_readRq, deq_fifo002);
    Module156 m156 <- mkModule156 (m135.cache_000_writeRs,
    m135.cache_000_removeVictim, m135.cache_000_getVictim,
    m28.transferUpDown000, m28.releaseDL000, m28.releaseUL000,
    m28.upLockGet000, m72.deq_fifo00031, m61.deq_fifo00021,
    m50.deq_fifo00011, m28.addRs000, m28.downLockGet000, m39.deq_fifo00001,
    m136.broadcast_parentChildren000, m28.registerDL000, m28.registerUL000,
    m135.cache_000_hasVictimSlot, m136.makeEnq_parentChildren000,
    m135.cache_000_writeRq, m28.downLockable000, m28.upLockable000,
    m135.cache_000_readRs, m71.deq_fifo00030, m60.deq_fifo00020,
    m49.deq_fifo00010, m38.deq_fifo00000, m28.downLockRssFull000,
    m135.cache_000_readRq, m31.deq_fifo0002);
    Module157 m157 <- mkModule157 (m137.cache_0000_writeRs,
    m137.cache_0000_removeVictim, m137.cache_0000_getVictim,
    m37.releaseUL0000, m137.cache_0000_writeRq, m37.upLockGet0000,
    m37.registerUL0000, m137.cache_0000_hasVictimSlot,
    m138.makeEnq_parentChildren0000, m37.downLockable0000,
    m37.upLockable0000, m137.cache_0000_readRs, m41.deq_fifo000000,
    m37.downLockRssFull0000, m137.cache_0000_readRq, m40.deq_fifo00002);

    Module158 m158 <- mkModule158 (m139.cache_0001_writeRs,
    m139.cache_0001_removeVictim, m139.cache_0001_getVictim,
    m48.releaseUL0001, m139.cache_0001_writeRq, m48.upLockGet0001,
    m48.registerUL0001, m139.cache_0001_hasVictimSlot,
    m140.makeEnq_parentChildren0001, m48.downLockable0001,
    m48.upLockable0001, m139.cache_0001_readRs, m52.deq_fifo000100,
    m48.downLockRssFull0001, m139.cache_0001_readRq, m51.deq_fifo00012);

    Module159 m159 <- mkModule159 (m141.cache_0002_writeRs,
    m141.cache_0002_removeVictim, m141.cache_0002_getVictim,
    m59.releaseUL0002, m141.cache_0002_writeRq, m59.upLockGet0002,
    m59.registerUL0002, m141.cache_0002_hasVictimSlot,
    m142.makeEnq_parentChildren0002, m59.downLockable0002,
    m59.upLockable0002, m141.cache_0002_readRs, m63.deq_fifo000200,
    m59.downLockRssFull0002, m141.cache_0002_readRq, m62.deq_fifo00022);

    Module160 m160 <- mkModule160 (m143.cache_0003_writeRs,
    m143.cache_0003_removeVictim, m143.cache_0003_getVictim,
    m70.releaseUL0003, m143.cache_0003_writeRq, m70.upLockGet0003,
    m70.registerUL0003, m143.cache_0003_hasVictimSlot,
    m144.makeEnq_parentChildren0003, m70.downLockable0003,
    m70.upLockable0003, m143.cache_0003_readRs, m74.deq_fifo000300,
    m70.downLockRssFull0003, m143.cache_0003_readRq, m73.deq_fifo00032);

    Module161 m161 <- mkModule161 (m145.cache_001_writeRs,
    m145.cache_001_removeVictim, m145.cache_001_getVictim,
    m85.transferUpDown001, m85.releaseDL001, m85.releaseUL001,
    m85.upLockGet001, m129.deq_fifo00131, m118.deq_fifo00121,
    m107.deq_fifo00111, m85.addRs001, m85.downLockGet001, m96.deq_fifo00101,
    m146.broadcast_parentChildren001, m85.registerDL001, m85.registerUL001,
    m145.cache_001_hasVictimSlot, m146.makeEnq_parentChildren001,
    m145.cache_001_writeRq, m85.downLockable001, m85.upLockable001,
    m145.cache_001_readRs, m128.deq_fifo00130, m117.deq_fifo00120,
    m106.deq_fifo00110, m95.deq_fifo00100, m85.downLockRssFull001,
    m145.cache_001_readRq, m88.deq_fifo0012);
    Module162 m162 <- mkModule162 (m147.cache_0010_writeRs,
    m147.cache_0010_removeVictim, m147.cache_0010_getVictim,
    m94.releaseUL0010, m147.cache_0010_writeRq, m94.upLockGet0010,
    m94.registerUL0010, m147.cache_0010_hasVictimSlot,
    m148.makeEnq_parentChildren0010, m94.downLockable0010,
    m94.upLockable0010, m147.cache_0010_readRs, m98.deq_fifo001000,
    m94.downLockRssFull0010, m147.cache_0010_readRq, m97.deq_fifo00102);

    Module163 m163 <- mkModule163 (m149.cache_0011_writeRs,
    m149.cache_0011_removeVictim, m149.cache_0011_getVictim,
    m105.releaseUL0011, m149.cache_0011_writeRq, m105.upLockGet0011,
    m105.registerUL0011, m149.cache_0011_hasVictimSlot,
    m150.makeEnq_parentChildren0011, m105.downLockable0011,
    m105.upLockable0011, m149.cache_0011_readRs, m109.deq_fifo001100,
    m105.downLockRssFull0011, m149.cache_0011_readRq, m108.deq_fifo00112);

    Module164 m164 <- mkModule164 (m151.cache_0012_writeRs,
    m151.cache_0012_removeVictim, m151.cache_0012_getVictim,
    m116.releaseUL0012, m151.cache_0012_writeRq, m116.upLockGet0012,
    m116.registerUL0012, m151.cache_0012_hasVictimSlot,
    m152.makeEnq_parentChildren0012, m116.downLockable0012,
    m116.upLockable0012, m151.cache_0012_readRs, m120.deq_fifo001200,
    m116.downLockRssFull0012, m151.cache_0012_readRq, m119.deq_fifo00122);

    Module165 m165 <- mkModule165 (m153.cache_0013_writeRs,
    m153.cache_0013_removeVictim, m153.cache_0013_getVictim,
    m127.releaseUL0013, m153.cache_0013_writeRq, m127.upLockGet0013,
    m127.registerUL0013, m153.cache_0013_hasVictimSlot,
    m154.makeEnq_parentChildren0013, m127.downLockable0013,
    m127.upLockable0013, m153.cache_0013_readRs, m131.deq_fifo001300,
    m127.downLockRssFull0013, m153.cache_0013_readRq, m130.deq_fifo00132);

        //// Initialization logic

    Reg#(Bool) init <- mkReg(False);

    Reg#(Bool) llInitDone <- mkReg(False);
    Reg#(Bit#(10)) llInitIndex <- mkReg(0);

    Reg#(Bool) l2InitDone0 <- mkReg(False);
    Reg#(Bit#(8)) l2InitIndex0 <- mkReg(0);
    Reg#(Bool) l2InitDone1 <- mkReg(False);
    Reg#(Bit#(8)) l2InitIndex1 <- mkReg(0);

    Reg#(Bool) l1InitDone0 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex0 <- mkReg(0);
    Reg#(Bool) l1InitDone1 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex1 <- mkReg(0);
    Reg#(Bool) l1InitDone2 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex2 <- mkReg(0);
    Reg#(Bool) l1InitDone3 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex3 <- mkReg(0);
    Reg#(Bool) l1InitDone4 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex4 <- mkReg(0);
    Reg#(Bool) l1InitDone5 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex5 <- mkReg(0);
    Reg#(Bool) l1InitDone6 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex6 <- mkReg(0);
    Reg#(Bool) l1InitDone7 <- mkReg(False);
    Reg#(Bit#(6)) l1InitIndex7 <- mkReg(0);

    function Struct22 llDefaultLine (Bit#(51) tagValue);
      return Struct22 { write: True,
                       addr: llInitIndex,
                       datain: Struct19 { tag: tagValue,
                                         value: Struct4 { mesi_owned: False,
                                                         mesi_status: 3'h1,
                                                         mesi_dir_st: 3'h1,
                                                         mesi_dir_sharers: 4'h0 }}};
    endfunction

    rule ll_info_do_init (!llInitDone);
        m1.putRq_infoRam_00_15 (llDefaultLine(15));
        m2.putRq_infoRam_00_14 (llDefaultLine(14));
        m3.putRq_infoRam_00_13 (llDefaultLine(13));
        m4.putRq_infoRam_00_12 (llDefaultLine(12));
        m5.putRq_infoRam_00_11 (llDefaultLine(11));
        m6.putRq_infoRam_00_10 (llDefaultLine(10));
        m7.putRq_infoRam_00_9 (llDefaultLine(9));
        m8.putRq_infoRam_00_8 (llDefaultLine(8));
        m9.putRq_infoRam_00_7 (llDefaultLine(7));
        m10.putRq_infoRam_00_6 (llDefaultLine(6));
        m11.putRq_infoRam_00_5 (llDefaultLine(5));
        m12.putRq_infoRam_00_4 (llDefaultLine(4));
        m13.putRq_infoRam_00_3 (llDefaultLine(3));
        m14.putRq_infoRam_00_2 (llDefaultLine(2));
        m15.putRq_infoRam_00_1 (llDefaultLine(1));
        m16.putRq_infoRam_00_0 (llDefaultLine(0));

        llInitIndex <= llInitIndex + 1;
        if (llInitIndex == 10'b1111111111) begin
            $display ("-- ll: initialization completed");
            llInitDone <= True;
        end
    endrule

    function Struct29 l2DefaultLine (Bit#(53) tagValue, Bit#(8) index);
      return Struct29 { write: True,
                       addr: index,
                       datain: Struct26 { tag: tagValue,
                                         value: Struct4 { mesi_owned: False,
                                                         mesi_status: 3'h1,
                                                         mesi_dir_st: 3'h1,
                                                         mesi_dir_sharers: 4'h0 }}};
    endfunction

    rule l2_info_do_init_0 (!l2InitDone0);
        m19.putRq_infoRam_000_7 (l2DefaultLine(7, l2InitIndex0));
        m20.putRq_infoRam_000_6 (l2DefaultLine(6, l2InitIndex0));
        m21.putRq_infoRam_000_5 (l2DefaultLine(5, l2InitIndex0));
        m22.putRq_infoRam_000_4 (l2DefaultLine(4, l2InitIndex0));
        m23.putRq_infoRam_000_3 (l2DefaultLine(3, l2InitIndex0));
        m24.putRq_infoRam_000_2 (l2DefaultLine(2, l2InitIndex0));
        m25.putRq_infoRam_000_1 (l2DefaultLine(1, l2InitIndex0));
        m26.putRq_infoRam_000_0 (l2DefaultLine(0, l2InitIndex0));

        l2InitIndex0 <= l2InitIndex0 + 1;
        if (l2InitIndex0 == 8'b11111111) begin
            $display ("-- l2_0: initialization completed");
            l2InitDone0 <= True;
        end
    endrule

    rule l2_info_do_init_1 (!l2InitDone1);
        m76.putRq_infoRam_001_7 (l2DefaultLine(7, l2InitIndex1));
        m77.putRq_infoRam_001_6 (l2DefaultLine(6, l2InitIndex1));
        m78.putRq_infoRam_001_5 (l2DefaultLine(5, l2InitIndex1));
        m79.putRq_infoRam_001_4 (l2DefaultLine(4, l2InitIndex1));
        m80.putRq_infoRam_001_3 (l2DefaultLine(3, l2InitIndex1));
        m81.putRq_infoRam_001_2 (l2DefaultLine(2, l2InitIndex1));
        m82.putRq_infoRam_001_1 (l2DefaultLine(1, l2InitIndex1));
        m83.putRq_infoRam_001_0 (l2DefaultLine(0, l2InitIndex1));

        l2InitIndex1 <= l2InitIndex1 + 1;
        if (l2InitIndex1 == 8'b11111111) begin
            $display ("-- l2_1: initialization completed");
            l2InitDone1 <= True;
        end
    endrule

    function Struct36 l1DefaultLine (Bit#(55) tagValue, Bit#(6) index);
      return Struct36 { write: True,
                       addr: index,
                       datain: Struct33 { tag: tagValue,
                                         value: Struct4 { mesi_owned: False,
                                                         mesi_status: 3'h1,
                                                         mesi_dir_st: 3'h1,
                                                         mesi_dir_sharers: 4'h0 }}};
    endfunction

    rule l1_info_do_init_0 (!l1InitDone0);
        m32.putRq_infoRam_0000_3 (l1DefaultLine(3, l1InitIndex0));
        m33.putRq_infoRam_0000_2 (l1DefaultLine(2, l1InitIndex0));
        m34.putRq_infoRam_0000_1 (l1DefaultLine(1, l1InitIndex0));
        m35.putRq_infoRam_0000_0 (l1DefaultLine(0, l1InitIndex0));
        l1InitIndex0 <= l1InitIndex0 + 1;
        if (l1InitIndex0 == 6'b111111) begin
            $display ("-- l1_0: initialization completed");
            l1InitDone0 <= True;
        end
    endrule

    rule l1_info_do_init_1 (!l1InitDone1);
        m43.putRq_infoRam_0001_3 (l1DefaultLine(3, l1InitIndex1));
        m44.putRq_infoRam_0001_2 (l1DefaultLine(2, l1InitIndex1));
        m45.putRq_infoRam_0001_1 (l1DefaultLine(1, l1InitIndex1));
        m46.putRq_infoRam_0001_0 (l1DefaultLine(0, l1InitIndex1));
        l1InitIndex1 <= l1InitIndex1 + 1;
        if (l1InitIndex1 == 6'b111111) begin
            $display ("-- l1_1: initialization completed");
            l1InitDone1 <= True;
        end
    endrule

    rule l1_info_do_init_2 (!l1InitDone2);
        m54.putRq_infoRam_0002_3 (l1DefaultLine(3, l1InitIndex2));
        m55.putRq_infoRam_0002_2 (l1DefaultLine(2, l1InitIndex2));
        m56.putRq_infoRam_0002_1 (l1DefaultLine(1, l1InitIndex2));
        m57.putRq_infoRam_0002_0 (l1DefaultLine(0, l1InitIndex2));
        l1InitIndex2 <= l1InitIndex1 + 1;
        if (l1InitIndex2 == 6'b111111) begin
            $display ("-- l1_2: initialization completed");
            l1InitDone2 <= True;
        end
    endrule

    rule l1_info_do_init_3 (!l1InitDone3);
        m65.putRq_infoRam_0003_3 (l1DefaultLine(3, l1InitIndex3));
        m66.putRq_infoRam_0003_2 (l1DefaultLine(2, l1InitIndex3));
        m67.putRq_infoRam_0003_1 (l1DefaultLine(1, l1InitIndex3));
        m68.putRq_infoRam_0003_0 (l1DefaultLine(0, l1InitIndex3));
        l1InitIndex3 <= l1InitIndex1 + 1;
        if (l1InitIndex3 == 6'b111111) begin
            $display ("-- l1_3: initialization completed");
            l1InitDone3 <= True;
        end
    endrule

    rule l1_info_do_init_4 (!l1InitDone4);
        m89.putRq_infoRam_0010_3 (l1DefaultLine(3, l1InitIndex4));
        m90.putRq_infoRam_0010_2 (l1DefaultLine(2, l1InitIndex4));
        m91.putRq_infoRam_0010_1 (l1DefaultLine(1, l1InitIndex4));
        m92.putRq_infoRam_0010_0 (l1DefaultLine(0, l1InitIndex4));
        l1InitIndex4 <= l1InitIndex4 + 1;
        if (l1InitIndex4 == 6'b111111) begin
            $display ("-- l1_4: initialization completed");
            l1InitDone4 <= True;
        end
    endrule

    rule l1_info_do_init_5 (!l1InitDone5);
        m100.putRq_infoRam_0011_3 (l1DefaultLine(3, l1InitIndex5));
        m101.putRq_infoRam_0011_2 (l1DefaultLine(2, l1InitIndex5));
        m102.putRq_infoRam_0011_1 (l1DefaultLine(1, l1InitIndex5));
        m103.putRq_infoRam_0011_0 (l1DefaultLine(0, l1InitIndex5));
        l1InitIndex5 <= l1InitIndex5 + 1;
        if (l1InitIndex5 == 6'b111111) begin
            $display ("-- l1_5: initialization completed");
            l1InitDone5 <= True;
        end
    endrule

    rule l1_info_do_init_6 (!l1InitDone6);
        m111.putRq_infoRam_0012_3 (l1DefaultLine(3, l1InitIndex6));
        m112.putRq_infoRam_0012_2 (l1DefaultLine(2, l1InitIndex6));
        m113.putRq_infoRam_0012_1 (l1DefaultLine(1, l1InitIndex6));
        m114.putRq_infoRam_0012_0 (l1DefaultLine(0, l1InitIndex6));
        l1InitIndex6 <= l1InitIndex6 + 1;
        if (l1InitIndex6 == 6'b111111) begin
            $display ("-- l1_6: initialization completed");
            l1InitDone6 <= True;
        end
    endrule

    rule l1_info_do_init_7 (!l1InitDone7);
        m122.putRq_infoRam_0013_3 (l1DefaultLine(3, l1InitIndex7));
        m123.putRq_infoRam_0013_2 (l1DefaultLine(2, l1InitIndex7));
        m124.putRq_infoRam_0013_1 (l1DefaultLine(1, l1InitIndex7));
        m125.putRq_infoRam_0013_0 (l1DefaultLine(0, l1InitIndex7));
        l1InitIndex7 <= l1InitIndex7 + 1;
        if (l1InitIndex7 == 6'b111111) begin
            $display ("-- l1_7: initialization completed");
            l1InitDone7 <= True;
        end
    endrule

    rule init_done (!init && llInitDone &&
                    l2InitDone0 && l2InitDone1 &&
                    l1InitDone0 && l1InitDone1 && l1InitDone2 && l1InitDone3 &&
                    l1InitDone4 && l1InitDone5 && l1InitDone6 && l1InitDone7);
        $display ("-- ALL: initialization completed");
        init <= True;
    endrule

    method Bool isInit ();
        return init;
    endmethod

    //// Interface
    method mem_enq_rq_0 = m41.enq_fifo000000;
    method mem_deq_rs_0 = m42.deq_fifo000002;
    method mem_enq_rq_1 = m52.enq_fifo000100;
    method mem_deq_rs_1 = m53.deq_fifo000102;
    method mem_enq_rq_2 = m63.enq_fifo000200;
    method mem_deq_rs_2 = m64.deq_fifo000202;
    method mem_enq_rq_3 = m74.enq_fifo000300;
    method mem_deq_rs_3 = m75.deq_fifo000302;

    method mem_enq_rq_4 = m98.enq_fifo001000;
    method mem_deq_rs_4 = m99.deq_fifo001002;
    method mem_enq_rq_5 = m109.enq_fifo001100;
    method mem_deq_rs_5 = m110.deq_fifo001102;
    method mem_enq_rq_6 = m120.enq_fifo001200;
    method mem_deq_rs_6 = m121.deq_fifo001202;
    method mem_enq_rq_7 = m131.enq_fifo001300;
    method mem_deq_rs_7 = m132.deq_fifo001302;

endmodule
