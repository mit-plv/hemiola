import Vector::*;
import BuildVector::*;
import FIFO::*;
import FIFOF::*;

import CC::*;

typedef Struct2 CCMsg;
typedef Bit#(6) CCMsgId;
typedef Bit#(64) CCAddr;
typedef Bit#(64) CCValue;
