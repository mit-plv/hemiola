CCIfc4.bsv