CC_L1LL8.bsv