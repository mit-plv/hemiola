CCWrapper_L1L2LL.bsv