CCWrapper.bsv