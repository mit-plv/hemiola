import Vector::*;
import BuildVector::*;
import FIFO::*;
import FIFOF::*;
import RWBramCore::*;
import SpecialFIFOs::*;

typedef 4 L1Num;

interface MemRqRs;
    method Action mem_enq_rq (Struct2 rq);
    method ActionValue#(Struct2) mem_deq_rs ();
endinterface

interface DMA;
    method Action dma_putRq (Struct21 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) dma_getRs ();
endinterface

interface CC;
    interface Vector#(L1Num, MemRqRs) l1Ifc;
    interface DMA llDma;
    method Bool isInit ();
endinterface

typedef struct { Bool rl_valid; Bit#(2) rl_cmidx; Struct2 rl_msg; Bool rl_line_valid; Struct3 rl_line;  } Struct1 deriving(Eq, Bits);
typedef struct { Bit#(2) enq_type; Bit#(2) enq_ch_idx; Struct2 enq_msg;  } Struct10 deriving(Eq, Bits);
typedef struct { Bool r_ul_rsb; Struct2 r_ul_msg; Bit#(2) r_ul_rsbTo;  } Struct11 deriving(Eq, Bits);
typedef struct { Bool r_dl_rsb; Struct2 r_dl_msg; Bit#(4) r_dl_rss_from; Bit#(4) r_dl_rsbTo;  } Struct12 deriving(Eq, Bits);
typedef struct { Bit#(4) cs_inds; Struct2 cs_msg;  } Struct13 deriving(Eq, Bits);
typedef struct { Bit#(64) r_dl_addr; Bit#(2) r_dl_midx; Struct2 r_dl_msg;  } Struct14 deriving(Eq, Bits);
typedef struct { Bool valid; Struct9 data;  } Struct15 deriving(Eq, Bits);
typedef struct { Bit#(4) cidx; Struct2 msg;  } Struct16 deriving(Eq, Bits);
typedef struct { Bit#(64) r_dl_addr; Bit#(4) r_dl_rss_from;  } Struct17 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(2) victim_idx; Struct3 victim_line;  } Struct18 deriving(Eq, Bits);
typedef struct { Bit#(49) tag; Struct4 value;  } Struct19 deriving(Eq, Bits);
typedef struct { Bit#(6) id; Bool type_; Bit#(64) addr; Vector#(4, Bit#(64)) value;  } Struct2 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(4) tm_way; Struct4 tm_value;  } Struct20 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(14) addr; Vector#(4, Bit#(64)) datain;  } Struct21 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(10) addr; Struct19 datain;  } Struct22 deriving(Eq, Bits);
typedef struct { Bool rl_valid; Bit#(2) rl_cmidx; Struct2 rl_msg; Bool rl_line_valid; Struct24 rl_line;  } Struct23 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_hit; Bit#(2) info_way; Bool info_write; Struct4 info; Bool value_write; Vector#(4, Bit#(64)) value;  } Struct24 deriving(Eq, Bits);
typedef struct { Bool victim_valid; Bit#(2) victim_idx; Struct24 victim_line;  } Struct25 deriving(Eq, Bits);
typedef struct { Bit#(51) tag; Struct4 value;  } Struct26 deriving(Eq, Bits);
typedef struct { Bool tm_hit; Bit#(2) tm_way; Struct4 tm_value;  } Struct27 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(10) addr; Vector#(4, Bit#(64)) datain;  } Struct28 deriving(Eq, Bits);
typedef struct { Bool write; Bit#(8) addr; Struct26 datain;  } Struct29 deriving(Eq, Bits);
typedef struct { Bit#(64) addr; Bool info_hit; Bit#(4) info_way; Bool info_write; Struct4 info; Bool value_write; Vector#(4, Bit#(64)) value;  } Struct3 deriving(Eq, Bits);
typedef struct { Bool mesi_owned; Bit#(3) mesi_status; Bit#(3) mesi_dir_st; Bit#(4) mesi_dir_sharers;  } Struct4 deriving(Eq, Bits);
typedef struct { Bool wl_valid; Bool wl_write_rq;  } Struct5 deriving(Eq, Bits);
typedef struct { Bool valid; Struct7 data;  } Struct6 deriving(Eq, Bits);
typedef struct { Bool dl_valid; Bool dl_rsb; Struct2 dl_msg; Bit#(4) dl_rss_from; Bit#(4) dl_rss_recv; Vector#(4, Struct2) dl_rss; Bit#(4) dl_rsbTo;  } Struct7 deriving(Eq, Bits);
typedef struct { Bit#(3) dir_st; Bit#(2) dir_excl; Bit#(4) dir_sharers;  } Struct8 deriving(Eq, Bits);
typedef struct { Bool ul_valid; Bool ul_rsb; Struct2 ul_msg; Bit#(2) ul_rsbTo;  } Struct9 deriving(Eq, Bits);

interface Module1;
    method Action putRq_infoRam_00_15 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_15 ();

endinterface

module mkModule1 (Module1);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_15 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_15 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module2;
    method Action putRq_infoRam_00_14 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_14 ();

endinterface

module mkModule2 (Module2);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_14 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_14 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module3;
    method Action putRq_infoRam_00_13 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_13 ();

endinterface

module mkModule3 (Module3);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_13 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_13 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module4;
    method Action putRq_infoRam_00_12 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_12 ();

endinterface

module mkModule4 (Module4);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_12 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_12 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module5;
    method Action putRq_infoRam_00_11 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_11 ();

endinterface

module mkModule5 (Module5);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_11 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_11 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module6;
    method Action putRq_infoRam_00_10 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_10 ();

endinterface

module mkModule6 (Module6);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_10 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_10 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module7;
    method Action putRq_infoRam_00_9 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_9 ();

endinterface

module mkModule7 (Module7);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_9 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_9 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module8;
    method Action putRq_infoRam_00_8 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_8 ();

endinterface

module mkModule8 (Module8);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_8 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_8 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module9;
    method Action putRq_infoRam_00_7 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_7 ();

endinterface

module mkModule9 (Module9);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_7 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_7 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module10;
    method Action putRq_infoRam_00_6 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_6 ();

endinterface

module mkModule10 (Module10);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_6 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_6 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module11;
    method Action putRq_infoRam_00_5 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_5 ();

endinterface

module mkModule11 (Module11);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_5 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_5 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module12;
    method Action putRq_infoRam_00_4 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_4 ();

endinterface

module mkModule12 (Module12);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_4 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_4 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module13;
    method Action putRq_infoRam_00_3 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_3 ();

endinterface

module mkModule13 (Module13);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_3 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module14;
    method Action putRq_infoRam_00_2 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_2 ();

endinterface

module mkModule14 (Module14);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_2 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module15;
    method Action putRq_infoRam_00_1 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_1 ();

endinterface

module mkModule15 (Module15);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_1 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module16;
    method Action putRq_infoRam_00_0 (Struct22 x_0);
    method ActionValue#(Struct19) getRs_infoRam_00_0 ();

endinterface

module mkModule16 (Module16);
    RWBramCore#(Bit#(10), Struct19) bram <- mkRWBramCore();

    method Action putRq_infoRam_00_0 (Struct22 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct19) getRs_infoRam_00_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module17;
    method Action putRq_dataRam_00 (Struct21 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_00 ();

endinterface

module mkModule17 (Module17);
    RWBramCore#(Bit#(14), Vector#(4, Bit#(64))) bram <- mkRWBramCore();

    method Action putRq_dataRam_00 (Struct21 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end

    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_00 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module18;
    method ActionValue#(Bool) upLockable00 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable00 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet00 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet00 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull00 ();
    method Action registerUL00 (Struct11 x_0);
    method Action releaseUL00 (Bit#(64) x_0);
    method Action registerDL00 (Struct12 x_0);
    method Action releaseDL00 (Bit#(64) x_0);
    method Action transferUpDown00 (Struct17 x_0);
    method Action addRs00 (Struct14 x_0);

endinterface

module mkModule18 (Module18);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable00 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable00 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).dl_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet00 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet00 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull00 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h2)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h2)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        ((((x_1)[(Bit#(2))'(2'h3)]).dl_rss_recv) ==
        (((x_1)[(Bit#(2))'(2'h3)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))))))));

        return x_2;
    endmethod

    method Action registerUL00 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL00 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL00 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).dl_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).dl_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).dl_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).dl_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL00 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown00 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(2) x_6 = ((! (((x_5)[(Bit#(2))'(2'h0)]).dl_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_5)[(Bit#(2))'(2'h1)]).dl_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_5)[(Bit#(2))'(2'h2)]).dl_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_5)[(Bit#(2))'(2'h3)]).dl_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs00 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct6 x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module19;
    method Action putRq_infoRam_000_3 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_3 ();

endinterface

module mkModule19 (Module19);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_3 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module20;
    method Action putRq_infoRam_000_2 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_2 ();

endinterface

module mkModule20 (Module20);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_2 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module21;
    method Action putRq_infoRam_000_1 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_1 ();

endinterface

module mkModule21 (Module21);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_1 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module22;
    method Action putRq_infoRam_000_0 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_000_0 ();

endinterface

module mkModule22 (Module22);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_000_0 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_000_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module23;
    method Action putRq_dataRam_000 (Struct28 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_000 ();

endinterface

module mkModule23 (Module23);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();

    method Action putRq_dataRam_000 (Struct28 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end

    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_000 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module24;
    method ActionValue#(Bool) upLockable000 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable000 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet000 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet000 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull000 ();
    method Action registerUL000 (Struct11 x_0);
    method Action releaseUL000 (Bit#(64) x_0);
    method Action registerDL000 (Struct12 x_0);
    method Action releaseDL000 (Bit#(64) x_0);
    method Action transferUpDown000 (Struct17 x_0);
    method Action addRs000 (Struct14 x_0);

endinterface

module mkModule24 (Module24);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable000 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable000 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet000 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet000 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull000 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL000 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL000 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL000 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL000 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown000 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs000 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module25;
    method Action enq_fifo0000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0000 ();

endinterface

module mkModule25 (Module25);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0000 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0000 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module26;
    method Action enq_fifo0001 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0001 ();

endinterface

module mkModule26 (Module26);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0001 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0001 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module27;
    method Action enq_fifo0002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0002 ();

endinterface

module mkModule27 (Module27);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0002 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0002 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module28;
    method Action enq_fifo00000 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00000 ();

endinterface

module mkModule28 (Module28);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00000 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00000 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module29;
    method Action enq_fifo00002 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00002 ();

endinterface

module mkModule29 (Module29);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00002 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00002 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module30;
    method Action putRq_infoRam_001_3 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_3 ();

endinterface

module mkModule30 (Module30);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_3 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module31;
    method Action putRq_infoRam_001_2 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_2 ();

endinterface

module mkModule31 (Module31);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_2 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module32;
    method Action putRq_infoRam_001_1 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_1 ();

endinterface

module mkModule32 (Module32);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_1 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module33;
    method Action putRq_infoRam_001_0 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_001_0 ();

endinterface

module mkModule33 (Module33);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_001_0 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_001_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module34;
    method Action putRq_dataRam_001 (Struct28 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_001 ();

endinterface

module mkModule34 (Module34);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();

    method Action putRq_dataRam_001 (Struct28 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end

    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_001 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module35;
    method ActionValue#(Bool) upLockable001 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable001 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet001 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet001 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull001 ();
    method Action registerUL001 (Struct11 x_0);
    method Action releaseUL001 (Bit#(64) x_0);
    method Action registerDL001 (Struct12 x_0);
    method Action releaseDL001 (Bit#(64) x_0);
    method Action transferUpDown001 (Struct17 x_0);
    method Action addRs001 (Struct14 x_0);

endinterface

module mkModule35 (Module35);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable001 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable001 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet001 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet001 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull001 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL001 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL001 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL001 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL001 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown001 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs001 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module36;
    method Action enq_fifo0010 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0010 ();

endinterface

module mkModule36 (Module36);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0010 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0010 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module37;
    method Action enq_fifo0011 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0011 ();

endinterface

module mkModule37 (Module37);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0011 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0011 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module38;
    method Action enq_fifo0012 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0012 ();

endinterface

module mkModule38 (Module38);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0012 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0012 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module39;
    method Action enq_fifo00100 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00100 ();

endinterface

module mkModule39 (Module39);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00100 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00100 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module40;
    method Action enq_fifo00102 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00102 ();

endinterface

module mkModule40 (Module40);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00102 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00102 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module41;
    method Action putRq_infoRam_002_3 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_002_3 ();

endinterface

module mkModule41 (Module41);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_002_3 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_002_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module42;
    method Action putRq_infoRam_002_2 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_002_2 ();

endinterface

module mkModule42 (Module42);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_002_2 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_002_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module43;
    method Action putRq_infoRam_002_1 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_002_1 ();

endinterface

module mkModule43 (Module43);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_002_1 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_002_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module44;
    method Action putRq_infoRam_002_0 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_002_0 ();

endinterface

module mkModule44 (Module44);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_002_0 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_002_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module45;
    method Action putRq_dataRam_002 (Struct28 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_002 ();

endinterface

module mkModule45 (Module45);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();

    method Action putRq_dataRam_002 (Struct28 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end

    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_002 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module46;
    method ActionValue#(Bool) upLockable002 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable002 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet002 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet002 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull002 ();
    method Action registerUL002 (Struct11 x_0);
    method Action releaseUL002 (Bit#(64) x_0);
    method Action registerDL002 (Struct12 x_0);
    method Action releaseDL002 (Bit#(64) x_0);
    method Action transferUpDown002 (Struct17 x_0);
    method Action addRs002 (Struct14 x_0);

endinterface

module mkModule46 (Module46);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable002 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable002 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet002 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet002 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull002 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL002 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL002 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL002 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL002 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown002 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs002 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module47;
    method Action enq_fifo0020 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0020 ();

endinterface

module mkModule47 (Module47);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0020 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0020 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module48;
    method Action enq_fifo0021 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0021 ();

endinterface

module mkModule48 (Module48);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0021 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0021 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module49;
    method Action enq_fifo0022 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0022 ();

endinterface

module mkModule49 (Module49);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0022 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0022 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module50;
    method Action enq_fifo00200 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00200 ();

endinterface

module mkModule50 (Module50);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00200 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00200 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module51;
    method Action enq_fifo00202 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00202 ();

endinterface

module mkModule51 (Module51);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00202 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00202 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module52;
    method Action putRq_infoRam_003_3 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_003_3 ();

endinterface

module mkModule52 (Module52);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_003_3 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_003_3 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module53;
    method Action putRq_infoRam_003_2 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_003_2 ();

endinterface

module mkModule53 (Module53);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_003_2 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_003_2 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module54;
    method Action putRq_infoRam_003_1 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_003_1 ();

endinterface

module mkModule54 (Module54);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_003_1 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_003_1 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module55;
    method Action putRq_infoRam_003_0 (Struct29 x_0);
    method ActionValue#(Struct26) getRs_infoRam_003_0 ();

endinterface

module mkModule55 (Module55);
    RWBramCore#(Bit#(8), Struct26) bram <- mkRWBramCore();

    method Action putRq_infoRam_003_0 (Struct29 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end
    endmethod

    method ActionValue#(Struct26) getRs_infoRam_003_0 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module56;
    method Action putRq_dataRam_003 (Struct28 x_0);
    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_003 ();

endinterface

module mkModule56 (Module56);
    RWBramCore#(Bit#(10), Vector#(4, Bit#(64))) bram <- mkRWBramCore();

    method Action putRq_dataRam_003 (Struct28 x_0);

        if (x_0.write) begin
        bram.wrReq(x_0.addr, x_0.datain);
        end else begin
        bram.rdReq(x_0.addr);

        end

    endmethod

    method ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_003 ();
    bram.deqRdResp ();
    let data = bram.rdResp ();
    return data;
    endmethod

endmodule

interface Module57;
    method ActionValue#(Bool) upLockable003 (Bit#(64) x_0);
    method ActionValue#(Bool) downLockable003 (Bit#(64) x_0);
    method ActionValue#(Struct15) upLockGet003 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockGet003 (Bit#(64) x_0);
    method ActionValue#(Struct6) downLockRssFull003 ();
    method Action registerUL003 (Struct11 x_0);
    method Action releaseUL003 (Bit#(64) x_0);
    method Action registerDL003 (Struct12 x_0);
    method Action releaseDL003 (Bit#(64) x_0);
    method Action transferUpDown003 (Struct17 x_0);
    method Action addRs003 (Struct14 x_0);

endinterface

module mkModule57 (Module57);
    Reg#(Vector#(4, Struct9)) uls <- mkReg(unpack(0));
    Reg#(Vector#(2, Struct7)) dls <- mkReg(unpack(0));

    // No rules in this module

    method ActionValue#(Bool) upLockable003 (Bit#(64) x_0);
        let x_1 = (uls);
        Bool x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ? ((Bool)'(True)) : ((!
        (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))))))));
        Bool x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Bool) downLockable003 (Bit#(64) x_0);
        let x_1 = (dls);
        Bool x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ? ((Bool)'(True))
        : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ? ((Bool)'(True)) :
        ((Bool)'(False))))));
        Bool x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bool)'(False)) : ((Bool)'(True))))));
        return (x_2) && (x_3);
    endmethod

    method ActionValue#(Struct15) upLockGet003 (Bit#(64) x_0);
        let x_1 = (uls);
        Struct15 x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h0)]}) :
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h1)]}) :
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h2)]}) :
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ? (Struct15
        {valid : (Bool)'(True), data : (x_1)[(Bit#(2))'(2'h3)]}) :
        ((Struct15)'(Struct15 {valid: False, data: Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}}))))))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockGet003 (Bit#(64) x_0);
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ? (Struct6
        {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method ActionValue#(Struct6) downLockRssFull003 ();
        let x_1 = (dls);
        Struct6 x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h0)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h0)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        ((((x_1)[(Bit#(1))'(1'h1)]).dl_rss_recv) ==
        (((x_1)[(Bit#(1))'(1'h1)]).dl_rss_from)) ? (Struct6 {valid :
        (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        return x_2;
    endmethod

    method Action registerUL003 (Struct11 x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = ((! (((x_1)[(Bit#(2))'(2'h0)]).ul_valid) ?
        ((Bit#(2))'(2'h0)) : ((! (((x_1)[(Bit#(2))'(2'h1)]).ul_valid) ?
        ((Bit#(2))'(2'h1)) : ((! (((x_1)[(Bit#(2))'(2'h2)]).ul_valid) ?
        ((Bit#(2))'(2'h2)) : ((! (((x_1)[(Bit#(2))'(2'h3)]).ul_valid) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2, Struct9 {ul_valid : (Bool)'(True), ul_rsb :
        (x_0).r_ul_rsb, ul_msg : (x_0).r_ul_msg, ul_rsbTo :
        (x_0).r_ul_rsbTo});

    endmethod

    method Action releaseUL003 (Bit#(64) x_0);
        let x_1 = (uls);
        Bit#(2) x_2 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_0)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        uls <= update (x_1, x_2,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));


    endmethod

    method Action registerDL003 (Struct12 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = ((! (((x_1)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_1)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_0).r_dl_rsb, dl_msg : (x_0).r_dl_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : (x_0).r_dl_rsbTo});

    endmethod

    method Action releaseDL003 (Bit#(64) x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == (x_0)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        dls <= update (x_1, x_2,
        (Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));


    endmethod

    method Action transferUpDown003 (Struct17 x_0);
        let x_1 = (uls);
        Bit#(64) x_2 = ((x_0).r_dl_addr);
        Bit#(2) x_3 = (((((x_1)[(Bit#(2))'(2'h0)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h0)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h0)) : (((((x_1)[(Bit#(2))'(2'h1)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h1)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h1)) : (((((x_1)[(Bit#(2))'(2'h2)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h2)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h2)) : (((((x_1)[(Bit#(2))'(2'h3)]).ul_valid) &&
        (((((x_1)[(Bit#(2))'(2'h3)]).ul_msg).addr) == (x_2)) ?
        ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));
        Struct9 x_4 = ((x_1)[x_3]);
        let x_5 = (dls);
        Bit#(1) x_6 = ((! (((x_5)[(Bit#(1))'(1'h0)]).dl_valid) ?
        ((Bit#(1))'(1'h0)) : ((! (((x_5)[(Bit#(1))'(1'h1)]).dl_valid) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        uls <= update (x_1, x_3,
        (Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        dls <= update (x_5, x_6, Struct7 {dl_valid : (Bool)'(True), dl_rsb :
        (x_4).ul_rsb, dl_msg : (x_4).ul_msg, dl_rss_from :
        (x_0).r_dl_rss_from, dl_rss_recv : (Bit#(4))'(4'h0), dl_rss :
        (Vector#(4, Struct2))'(vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})),
        dl_rsbTo : {((Bit#(2))'(2'h2)),((x_4).ul_rsbTo)}});

    endmethod

    method Action addRs003 (Struct14 x_0);
        let x_1 = (dls);
        Bit#(1) x_2 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h0)) : (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        ((Bit#(1))'(1'h1)) : ((Bit#(1))'(1'h0))))));
        Struct6 x_3 = (((((x_1)[(Bit#(1))'(1'h0)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h0)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h0)]}) :
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_valid) &&
        (((((x_1)[(Bit#(1))'(1'h1)]).dl_msg).addr) == ((x_0).r_dl_addr)) ?
        (Struct6 {valid : (Bool)'(True), data : (x_1)[(Bit#(1))'(1'h1)]}) :
        ((Struct6)'(Struct6 {valid: False, data: Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}}))))));

        Struct7 x_4 = ((x_3).data);
        dls <= update (x_1, x_2, Struct7 {dl_valid : (x_4).dl_valid, dl_rsb :
        (x_4).dl_rsb, dl_msg : (x_4).dl_msg, dl_rss_from : (x_4).dl_rss_from,
        dl_rss_recv : ((x_4).dl_rss_recv) | (((Bit#(4))'(4'h1)) <<
        ((x_0).r_dl_midx)), dl_rss : update ((x_4).dl_rss, (x_0).r_dl_midx,
        (x_0).r_dl_msg), dl_rsbTo : (x_4).dl_rsbTo});

    endmethod

endmodule

interface Module58;
    method Action enq_fifo0030 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0030 ();

endinterface

module mkModule58 (Module58);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0030 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0030 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module59;
    method Action enq_fifo0031 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0031 ();

endinterface

module mkModule59 (Module59);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0031 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0031 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module60;
    method Action enq_fifo0032 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo0032 ();

endinterface

module mkModule60 (Module60);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo0032 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo0032 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module61;
    method Action enq_fifo00300 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00300 ();

endinterface

module mkModule61 (Module61);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00300 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00300 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module62;
    method Action enq_fifo00302 (Struct2 x_0);
    method ActionValue#(Struct2) deq_fifo00302 ();

endinterface

module mkModule62 (Module62);
    FIFOF#(Struct2) pff <- mkPipelineFIFOF();

    method Action enq_fifo00302 (Struct2 x_0);
    pff.enq(x_0);
    endmethod

    method ActionValue#(Struct2) deq_fifo00302 ();
    pff.deq();
    return pff.first();
    endmethod


endmodule

interface Module63;
    method Action cache_00_readRq (Bit#(64) x_0);
    method ActionValue#(Struct3) cache_00_readRs ();
    method Action cache_00_writeRq (Struct3 x_0);
    method ActionValue#(Struct3) cache_00_writeRs ();
    method ActionValue#(Bool) cache_00_hasVictimSlot ();
    method ActionValue#(Struct3) cache_00_getVictim ();
    method Action cache_00_removeVictim (Bit#(64) x_0);

endinterface


module mkModule63#(function Action putRq_infoRam_00_15(Struct22 _),
  function Action putRq_infoRam_00_14(Struct22 _),
  function Action putRq_infoRam_00_13(Struct22 _),
  function Action putRq_infoRam_00_12(Struct22 _),
  function Action putRq_infoRam_00_11(Struct22 _),
  function Action putRq_infoRam_00_10(Struct22 _),
  function Action putRq_infoRam_00_9(Struct22 _),
  function Action putRq_infoRam_00_8(Struct22 _),
  function Action putRq_infoRam_00_7(Struct22 _),
  function Action putRq_infoRam_00_6(Struct22 _),
  function Action putRq_infoRam_00_5(Struct22 _),
  function Action putRq_infoRam_00_4(Struct22 _),
  function Action putRq_infoRam_00_3(Struct22 _),
  function Action putRq_infoRam_00_2(Struct22 _),
  function Action putRq_infoRam_00_1(Struct22 _),
  function Action putRq_infoRam_00_0(Struct22 _),
  function ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_00(),
  function Action putRq_dataRam_00(Struct21 _),
  function ActionValue#(Struct19) getRs_infoRam_00_15(),
  function ActionValue#(Struct19) getRs_infoRam_00_14(),
  function ActionValue#(Struct19) getRs_infoRam_00_13(),
  function ActionValue#(Struct19) getRs_infoRam_00_12(),
  function ActionValue#(Struct19) getRs_infoRam_00_11(),
  function ActionValue#(Struct19) getRs_infoRam_00_10(),
  function ActionValue#(Struct19) getRs_infoRam_00_9(),
  function ActionValue#(Struct19) getRs_infoRam_00_8(),
  function ActionValue#(Struct19) getRs_infoRam_00_7(),
  function ActionValue#(Struct19) getRs_infoRam_00_6(),
  function ActionValue#(Struct19) getRs_infoRam_00_5(),
  function ActionValue#(Struct19) getRs_infoRam_00_4(),
  function ActionValue#(Struct19) getRs_infoRam_00_3(),
  function ActionValue#(Struct19) getRs_infoRam_00_2(),
  function ActionValue#(Struct19) getRs_infoRam_00_1(),
  function ActionValue#(Struct19) getRs_infoRam_00_0()) (Module63);
    Reg#(Bit#(2)) readStage_00 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_00 <- mkReg(unpack(0));
    Reg#(Struct3) readLine_00 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_00 <- mkReg(unpack(0));
    Reg#(Struct3) writeLine_00 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct18)) victims_00 <- mkReg(unpack(0));
    Reg#(Struct3) victimLine_00 <- mkReg(unpack(0));
    Reg#(Bit#(4)) victimWay_00 <- mkReg(unpack(0));

    rule read_tagmatch_00;
        let x_0 = (readStage_00);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_00);
        Bit#(49) x_2 = ((x_1)[63:15]);
        Bit#(10) x_3 = ((x_1)[14:5]);
        Vector#(16, Struct19) x_4 =
        ((Vector#(16, Struct19))'(vec(Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_00_0();
        Vector#(16, Struct19) x_6 = (update (x_4, (Bit#(4))'(4'h0), x_5));
        let x_7 <- getRs_infoRam_00_1();
        Vector#(16, Struct19) x_8 = (update (x_6, (Bit#(4))'(4'h1), x_7));
        let x_9 <- getRs_infoRam_00_2();
        Vector#(16, Struct19) x_10 = (update (x_8, (Bit#(4))'(4'h2), x_9));

        let x_11 <- getRs_infoRam_00_3();
        Vector#(16, Struct19) x_12 = (update (x_10, (Bit#(4))'(4'h3), x_11));

        let x_13 <- getRs_infoRam_00_4();
        Vector#(16, Struct19) x_14 = (update (x_12, (Bit#(4))'(4'h4), x_13));

        let x_15 <- getRs_infoRam_00_5();
        Vector#(16, Struct19) x_16 = (update (x_14, (Bit#(4))'(4'h5), x_15));

        let x_17 <- getRs_infoRam_00_6();
        Vector#(16, Struct19) x_18 = (update (x_16, (Bit#(4))'(4'h6), x_17));

        let x_19 <- getRs_infoRam_00_7();
        Vector#(16, Struct19) x_20 = (update (x_18, (Bit#(4))'(4'h7), x_19));

        let x_21 <- getRs_infoRam_00_8();
        Vector#(16, Struct19) x_22 = (update (x_20, (Bit#(4))'(4'h8), x_21));

        let x_23 <- getRs_infoRam_00_9();
        Vector#(16, Struct19) x_24 = (update (x_22, (Bit#(4))'(4'h9), x_23));

        let x_25 <- getRs_infoRam_00_10();
        Vector#(16, Struct19) x_26 = (update (x_24, (Bit#(4))'(4'ha), x_25));

        let x_27 <- getRs_infoRam_00_11();
        Vector#(16, Struct19) x_28 = (update (x_26, (Bit#(4))'(4'hb), x_27));

        let x_29 <- getRs_infoRam_00_12();
        Vector#(16, Struct19) x_30 = (update (x_28, (Bit#(4))'(4'hc), x_29));

        let x_31 <- getRs_infoRam_00_13();
        Vector#(16, Struct19) x_32 = (update (x_30, (Bit#(4))'(4'hd), x_31));

        let x_33 <- getRs_infoRam_00_14();
        Vector#(16, Struct19) x_34 = (update (x_32, (Bit#(4))'(4'he), x_33));

        let x_35 <- getRs_infoRam_00_15();
        Vector#(16, Struct19) x_36 = (update (x_34, (Bit#(4))'(4'hf), x_35));

        Struct20 x_37 = (((((x_36)[(Bit#(4))'(4'h0)]).tag) == (x_2) ?
        (Struct20 {tm_hit : (Bool)'(True), tm_way : (Bit#(4))'(4'h0),
        tm_value : ((x_36)[(Bit#(4))'(4'h0)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h1)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h1), tm_value :
        ((x_36)[(Bit#(4))'(4'h1)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h2)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h2), tm_value :
        ((x_36)[(Bit#(4))'(4'h2)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h3)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h3), tm_value :
        ((x_36)[(Bit#(4))'(4'h3)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h4)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h4), tm_value :
        ((x_36)[(Bit#(4))'(4'h4)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h5)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h5), tm_value :
        ((x_36)[(Bit#(4))'(4'h5)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h6)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h6), tm_value :
        ((x_36)[(Bit#(4))'(4'h6)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h7)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h7), tm_value :
        ((x_36)[(Bit#(4))'(4'h7)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h8)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h8), tm_value :
        ((x_36)[(Bit#(4))'(4'h8)]).value}) :
        (((((x_36)[(Bit#(4))'(4'h9)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'h9), tm_value :
        ((x_36)[(Bit#(4))'(4'h9)]).value}) :
        (((((x_36)[(Bit#(4))'(4'ha)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'ha), tm_value :
        ((x_36)[(Bit#(4))'(4'ha)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hb)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hb), tm_value :
        ((x_36)[(Bit#(4))'(4'hb)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hc)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hc), tm_value :
        ((x_36)[(Bit#(4))'(4'hc)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hd)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hd), tm_value :
        ((x_36)[(Bit#(4))'(4'hd)]).value}) :
        (((((x_36)[(Bit#(4))'(4'he)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'he), tm_value :
        ((x_36)[(Bit#(4))'(4'he)]).value}) :
        (((((x_36)[(Bit#(4))'(4'hf)]).tag) == (x_2) ? (Struct20 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(4))'(4'hf), tm_value :
        ((x_36)[(Bit#(4))'(4'hf)]).value}) :
        ((Struct20)'(Struct20 {tm_hit: False, tm_way: 4'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))))))))))))))))))))))))))));

        readLine_00 <= Struct3 {addr : x_1, info_hit : (x_37).tm_hit,
        info_way : (x_37).tm_way, info_write : (Bool)'(False), info :
        (x_37).tm_value, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        if ((x_37).tm_hit) begin

            readStage_00 <= (Bit#(2))'(2'h2);
            let x_38 <- putRq_dataRam_00(Struct21 {write : (Bool)'(False),
            addr : {(x_3),((x_37).tm_way)}, datain :
            (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

        end else begin
        readStage_00 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_00;
        let x_0 = (readStage_00);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_00 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_00();
        let x_2 = (readLine_00);
        readLine_00 <= Struct3 {addr : (x_2).addr, info_hit : (x_2).info_hit,
        info_way : (x_2).info_way, info_write : (x_2).info_write, info :
        (x_2).info, value_write : (Bool)'(False), value : x_1};

    endrule

    rule write_info_hit_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_00);
        when ((x_1).info_hit, noAction);
        writeStage_00 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(49) x_3 = ((x_2)[63:15]);
        Bit#(10) x_4 = ((x_2)[14:5]);
        Bit#(4) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct22 x_6 = (Struct22 {write : (Bool)'(True), addr : x_4,
            datain : Struct19 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(4))'(4'h0))) begin
            let x_7 <- putRq_infoRam_00_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h1))) begin
            let x_9 <- putRq_infoRam_00_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h2))) begin
            let x_11 <- putRq_infoRam_00_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h3))) begin
            let x_13 <- putRq_infoRam_00_3(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h4))) begin
            let x_15 <- putRq_infoRam_00_4(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h5))) begin
            let x_17 <- putRq_infoRam_00_5(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h6))) begin
            let x_19 <- putRq_infoRam_00_6(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h7))) begin
            let x_21 <- putRq_infoRam_00_7(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h8))) begin
            let x_23 <- putRq_infoRam_00_8(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h9))) begin
            let x_25 <- putRq_infoRam_00_9(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'ha))) begin
            let x_27 <- putRq_infoRam_00_10(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hb))) begin
            let x_29 <- putRq_infoRam_00_11(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hc))) begin
            let x_31 <- putRq_infoRam_00_12(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hd))) begin
            let x_33 <- putRq_infoRam_00_13(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'he))) begin
            let x_35 <- putRq_infoRam_00_14(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hf))) begin
            let x_37 <- putRq_infoRam_00_15(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_40 <- putRq_dataRam_00(Struct21 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_00);
        when (! ((x_1).info_hit), noAction);
        writeStage_00 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(10) x_3 = ((x_2)[14:5]);
        Struct22 x_4 = (Struct22 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct19)'(Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_00_0(x_4);
        let x_6 <- putRq_infoRam_00_1(x_4);
        let x_7 <- putRq_infoRam_00_2(x_4);
        let x_8 <- putRq_infoRam_00_3(x_4);
        let x_9 <- putRq_infoRam_00_4(x_4);
        let x_10 <- putRq_infoRam_00_5(x_4);
        let x_11 <- putRq_infoRam_00_6(x_4);
        let x_12 <- putRq_infoRam_00_7(x_4);
        let x_13 <- putRq_infoRam_00_8(x_4);
        let x_14 <- putRq_infoRam_00_9(x_4);
        let x_15 <- putRq_infoRam_00_10(x_4);
        let x_16 <- putRq_infoRam_00_11(x_4);
        let x_17 <- putRq_infoRam_00_12(x_4);
        let x_18 <- putRq_infoRam_00_13(x_4);
        let x_19 <- putRq_infoRam_00_14(x_4);
        let x_20 <- putRq_infoRam_00_15(x_4);

    endrule

    rule write_info_miss_rep_rs_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_00 <= (Bit#(3))'(3'h3);
        Vector#(16, Struct19) x_1 =
        ((Vector#(16, Struct19))'(vec(Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_00_0();
        Vector#(16, Struct19) x_3 = (update (x_1, (Bit#(4))'(4'h0), x_2));
        let x_4 <- getRs_infoRam_00_1();
        Vector#(16, Struct19) x_5 = (update (x_3, (Bit#(4))'(4'h1), x_4));
        let x_6 <- getRs_infoRam_00_2();
        Vector#(16, Struct19) x_7 = (update (x_5, (Bit#(4))'(4'h2), x_6));
        let x_8 <- getRs_infoRam_00_3();
        Vector#(16, Struct19) x_9 = (update (x_7, (Bit#(4))'(4'h3), x_8));
        let x_10 <- getRs_infoRam_00_4();
        Vector#(16, Struct19) x_11 = (update (x_9, (Bit#(4))'(4'h4), x_10));

        let x_12 <- getRs_infoRam_00_5();
        Vector#(16, Struct19) x_13 = (update (x_11, (Bit#(4))'(4'h5), x_12));

        let x_14 <- getRs_infoRam_00_6();
        Vector#(16, Struct19) x_15 = (update (x_13, (Bit#(4))'(4'h6), x_14));

        let x_16 <- getRs_infoRam_00_7();
        Vector#(16, Struct19) x_17 = (update (x_15, (Bit#(4))'(4'h7), x_16));

        let x_18 <- getRs_infoRam_00_8();
        Vector#(16, Struct19) x_19 = (update (x_17, (Bit#(4))'(4'h8), x_18));

        let x_20 <- getRs_infoRam_00_9();
        Vector#(16, Struct19) x_21 = (update (x_19, (Bit#(4))'(4'h9), x_20));

        let x_22 <- getRs_infoRam_00_10();
        Vector#(16, Struct19) x_23 = (update (x_21, (Bit#(4))'(4'ha), x_22));

        let x_24 <- getRs_infoRam_00_11();
        Vector#(16, Struct19) x_25 = (update (x_23, (Bit#(4))'(4'hb), x_24));

        let x_26 <- getRs_infoRam_00_12();
        Vector#(16, Struct19) x_27 = (update (x_25, (Bit#(4))'(4'hc), x_26));

        let x_28 <- getRs_infoRam_00_13();
        Vector#(16, Struct19) x_29 = (update (x_27, (Bit#(4))'(4'hd), x_28));

        let x_30 <- getRs_infoRam_00_14();
        Vector#(16, Struct19) x_31 = (update (x_29, (Bit#(4))'(4'he), x_30));

        let x_32 <- getRs_infoRam_00_15();
        Vector#(16, Struct19) x_33 = (update (x_31, (Bit#(4))'(4'hf), x_32));

        Bit#(4) x_34 = ((((((x_33)[(Bit#(4))'(4'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h0)) :
        ((((((x_33)[(Bit#(4))'(4'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h1)) :
        ((((((x_33)[(Bit#(4))'(4'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h2)) :
        ((((((x_33)[(Bit#(4))'(4'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h3)) :
        ((((((x_33)[(Bit#(4))'(4'h4)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h4)) :
        ((((((x_33)[(Bit#(4))'(4'h5)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h5)) :
        ((((((x_33)[(Bit#(4))'(4'h6)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h6)) :
        ((((((x_33)[(Bit#(4))'(4'h7)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h7)) :
        ((((((x_33)[(Bit#(4))'(4'h8)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h8)) :
        ((((((x_33)[(Bit#(4))'(4'h9)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'h9)) :
        ((((((x_33)[(Bit#(4))'(4'ha)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'ha)) :
        ((((((x_33)[(Bit#(4))'(4'hb)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hb)) :
        ((((((x_33)[(Bit#(4))'(4'hc)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hc)) :
        ((((((x_33)[(Bit#(4))'(4'hd)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hd)) :
        ((((((x_33)[(Bit#(4))'(4'he)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'he)) :
        ((((((x_33)[(Bit#(4))'(4'hf)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(4))'(4'hf)) :
        ((Bit#(4))'(4'h0))))))))))))))))))))))))))))))))));
        let x_35 = (writeLine_00);
        Bit#(64) x_36 = ((x_35).addr);
        Bit#(10) x_37 = ((x_36)[14:5]);
        Struct19 x_38 = ((x_33)[x_34]);
        Bit#(49) x_39 = ((x_38).tag);
        Struct4 x_40 = ((x_38).value);
        victimWay_00 <= x_34;
        victimLine_00 <= Struct3 {addr :
        {(x_39),({(x_37),((Bit#(5))'(5'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(4))'(4'h0), info_write : (Bool)'(False), info :
        x_40, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        let x_41 <- putRq_dataRam_00(Struct21 {write : (Bool)'(False), addr :
        {(x_37),(x_34)}, datain :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

    endrule

    rule write_victim_rs_00;
        let x_0 = (writeStage_00);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_00);
        writeStage_00 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(49) x_3 = ((x_2)[63:15]);
        Bit#(10) x_4 = ((x_2)[14:5]);
        let x_5 = (victimWay_00);
        let x_6 = (victims_00);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_00();
        let x_9 = (victimLine_00);
        victims_00 <= update (x_6, x_7, Struct18 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct3 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_00 <= Struct3 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct22 x_10 = (Struct22 {write : (Bool)'(True), addr : x_4,
            datain : Struct19 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(4))'(4'h0))) begin
            let x_11 <- putRq_infoRam_00_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h1))) begin
            let x_13 <- putRq_infoRam_00_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h2))) begin
            let x_15 <- putRq_infoRam_00_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h3))) begin
            let x_17 <- putRq_infoRam_00_3(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h4))) begin
            let x_19 <- putRq_infoRam_00_4(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h5))) begin
            let x_21 <- putRq_infoRam_00_5(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h6))) begin
            let x_23 <- putRq_infoRam_00_6(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h7))) begin
            let x_25 <- putRq_infoRam_00_7(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h8))) begin
            let x_27 <- putRq_infoRam_00_8(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'h9))) begin
            let x_29 <- putRq_infoRam_00_9(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'ha))) begin
            let x_31 <- putRq_infoRam_00_10(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hb))) begin
            let x_33 <- putRq_infoRam_00_11(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hc))) begin
            let x_35 <- putRq_infoRam_00_12(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hd))) begin
            let x_37 <- putRq_infoRam_00_13(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'he))) begin
            let x_39 <- putRq_infoRam_00_14(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(4))'(4'hf))) begin
            let x_41 <- putRq_infoRam_00_15(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_44 <- putRq_dataRam_00(Struct21 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_00_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_00);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_00);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_00);
        Struct18 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_00 <= (Bit#(2))'(2'h3);
        readLine_00 <= (x_4).victim_line;

        end else begin

            Struct18 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_00 <= (Bit#(2))'(2'h3);
                readLine_00 <= (x_5).victim_line;

            end else begin

                Struct18 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_00 <= (Bit#(2))'(2'h3);
                    readLine_00 <= (x_6).victim_line;

                end else begin

                    Struct18 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_00 <= (Bit#(2))'(2'h3);
                        readLine_00 <= (x_7).victim_line;

                    end else begin

                        readStage_00 <= (Bit#(2))'(2'h1);
                        readAddr_00 <= x_0;
                        Bit#(10) x_8 = ((x_0)[14:5]);
                        Struct22 x_9 = (Struct22 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct19)'(Struct19 {tag: 49'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_00_0(x_9);
                        let x_11 <- putRq_infoRam_00_1(x_9);
                        let x_12 <- putRq_infoRam_00_2(x_9);
                        let x_13 <- putRq_infoRam_00_3(x_9);
                        let x_14 <- putRq_infoRam_00_4(x_9);
                        let x_15 <- putRq_infoRam_00_5(x_9);
                        let x_16 <- putRq_infoRam_00_6(x_9);
                        let x_17 <- putRq_infoRam_00_7(x_9);
                        let x_18 <- putRq_infoRam_00_8(x_9);
                        let x_19 <- putRq_infoRam_00_9(x_9);
                        let x_20 <- putRq_infoRam_00_10(x_9);
                        let x_21 <- putRq_infoRam_00_11(x_9);
                        let x_22 <- putRq_infoRam_00_12(x_9);
                        let x_23 <- putRq_infoRam_00_13(x_9);
                        let x_24 <- putRq_infoRam_00_14(x_9);
                        let x_25 <- putRq_infoRam_00_15(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct3) cache_00_readRs ();
        let x_1 = (readStage_00);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_00 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_00);
        return x_2;
    endmethod

    method Action cache_00_writeRq (Struct3 x_0);
        let x_1 = (readStage_00);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_00);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_00);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct18 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct3 x_6 = (Struct3 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) : ((Bit#(3))'(3'h1)));

            writeLine_00 <= x_6;
            victims_00 <= update (x_3, (Bit#(2))'(2'h0), Struct18
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct18 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct3 x_8 = (Struct3 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_00 <= x_8;
                victims_00 <= update (x_3, (Bit#(2))'(2'h1), Struct18
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct18 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct3 x_10 = (Struct3 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_00 <= x_10;
                    victims_00 <= update (x_3, (Bit#(2))'(2'h2), Struct18
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct18 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct3 x_12 = (Struct3 {addr : (x_0).addr, info_hit
                        : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_00 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_00 <= x_12;
                        victims_00 <= update (x_3, (Bit#(2))'(2'h3), Struct18
                        {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h3),
                        victim_line : x_12});

                    end else begin
                    writeStage_00 <= (Bit#(3))'(3'h1);
                    writeLine_00 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct3) cache_00_writeRs ();
        let x_1 = (writeStage_00);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_00 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_00);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_00_hasVictimSlot ();
        let x_1 = (victims_00);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct3) cache_00_getVictim ();
        let x_1 = (victims_00);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct3 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_00_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_00);
        Struct18 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_00 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct18)'(Struct18 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


        end else begin

            Struct18 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_00 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct18)'(Struct18 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


            end else begin

                Struct18 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_00 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct18)'(Struct18 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                end else begin

                    Struct18 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_00 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct18)'(Struct18 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module64;
    method Action makeEnq_parentChildren00 (Struct10 x_0);
    method Action broadcast_parentChildren00 (Struct13 x_0);

endinterface


module mkModule64#(function Action enq_fifo0002(Struct2 _),
  function Action enq_fifo0012(Struct2 _),
  function Action enq_fifo0022(Struct2 _),
  function Action enq_fifo0032(Struct2 _),
  function Action enq_fifo001(Struct2 _),
  function Action enq_fifo000(Struct2 _)) (Module64);

    // No rules in this module

    method Action makeEnq_parentChildren00 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo000((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo001((x_0).enq_msg);

            end else begin

                Bit#(2) x_3 = ((x_0).enq_ch_idx);
                Struct2 x_4 = ((x_0).enq_msg);
                if ((x_3) == ((Bit#(2))'(2'h3))) begin
                let x_5 <- enq_fifo0032(x_4);

                end else begin

                    if ((x_3) == ((Bit#(2))'(2'h2))) begin
                    let x_6 <- enq_fifo0022(x_4);

                    end else begin

                        if ((x_3) == ((Bit#(2))'(2'h1))) begin
                        let x_7 <- enq_fifo0012(x_4);

                        end else begin

                            if ((x_3) == ((Bit#(2))'(2'h0))) begin
                            let x_8 <- enq_fifo0002(x_4);

                            end else begin

                            end

                        end

                    end

                end

            end

        end

    endmethod

    method Action broadcast_parentChildren00 (Struct13 x_0);
        Bit#(4) x_1 = ((x_0).cs_inds);
        Struct2 x_2 = ((x_0).cs_msg);
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == (x_1))
        begin
        let x_3 <- enq_fifo0032(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == (x_1))
        begin
        let x_5 <- enq_fifo0022(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == (x_1))
        begin
        let x_7 <- enq_fifo0012(x_2);

        end else begin

        end
        if (((x_1) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == (x_1))
        begin
        let x_9 <- enq_fifo0002(x_2);

        end else begin

        end

    endmethod

endmodule

interface Module65;
    method Action cache_000_readRq (Bit#(64) x_0);
    method ActionValue#(Struct24) cache_000_readRs ();
    method Action cache_000_writeRq (Struct24 x_0);
    method ActionValue#(Struct24) cache_000_writeRs ();
    method ActionValue#(Bool) cache_000_hasVictimSlot ();
    method ActionValue#(Struct24) cache_000_getVictim ();
    method Action cache_000_removeVictim (Bit#(64) x_0);

endinterface


module mkModule65#(function Action putRq_infoRam_000_3(Struct29 _),
  function Action putRq_infoRam_000_2(Struct29 _),
  function Action putRq_infoRam_000_1(Struct29 _),
  function Action putRq_infoRam_000_0(Struct29 _),
  function ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_000(),
  function Action putRq_dataRam_000(Struct28 _),
  function ActionValue#(Struct26) getRs_infoRam_000_3(),
  function ActionValue#(Struct26) getRs_infoRam_000_2(),
  function ActionValue#(Struct26) getRs_infoRam_000_1(),
  function ActionValue#(Struct26) getRs_infoRam_000_0()) (Module65);
    Reg#(Bit#(2)) readStage_000 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_000 <- mkReg(unpack(0));
    Reg#(Struct24) readLine_000 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_000 <- mkReg(unpack(0));
    Reg#(Struct24) writeLine_000 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct25)) victims_000 <- mkReg(unpack(0));
    Reg#(Struct24) victimLine_000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_000 <- mkReg(unpack(0));

    rule read_tagmatch_000;
        let x_0 = (readStage_000);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_000);
        Bit#(51) x_2 = ((x_1)[63:13]);
        Bit#(8) x_3 = ((x_1)[12:5]);
        Vector#(4, Struct26) x_4 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_000_0();
        Vector#(4, Struct26) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_000_1();
        Vector#(4, Struct26) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_000_2();
        Vector#(4, Struct26) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_000_3();
        Vector#(4, Struct26) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct27 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct27 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct27)'(Struct27 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_000 <= Struct24 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        if ((x_13).tm_hit) begin

            readStage_000 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_000(Struct28 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain :
            (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

        end else begin
        readStage_000 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_000;
        let x_0 = (readStage_000);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_000 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_000();
        let x_2 = (readLine_000);
        readLine_000 <= Struct24 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_000);
        when ((x_1).info_hit, noAction);
        writeStage_000 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct29 x_6 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_000_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_000_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_000_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_000_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_000(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_000);
        when (! ((x_1).info_hit), noAction);
        writeStage_000 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Struct29 x_4 = (Struct29 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_000_0(x_4);
        let x_6 <- putRq_infoRam_000_1(x_4);
        let x_7 <- putRq_infoRam_000_2(x_4);
        let x_8 <- putRq_infoRam_000_3(x_4);

    endrule

    rule write_info_miss_rep_rs_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_000 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct26) x_1 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_000_0();
        Vector#(4, Struct26) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_000_1();
        Vector#(4, Struct26) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_000_2();
        Vector#(4, Struct26) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_000_3();
        Vector#(4, Struct26) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_000);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(8) x_13 = ((x_12)[12:5]);
        Struct26 x_14 = ((x_9)[x_10]);
        Bit#(51) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_000 <= x_10;
        victimLine_000 <= Struct24 {addr :
        {(x_15),({(x_13),((Bit#(5))'(5'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        let x_17 <- putRq_dataRam_000(Struct28 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

    endrule

    rule write_victim_rs_000;
        let x_0 = (writeStage_000);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_000);
        writeStage_000 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        let x_5 = (victimWay_000);
        let x_6 = (victims_000);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_000();
        let x_9 = (victimLine_000);
        victims_000 <= update (x_6, x_7, Struct25 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct24 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_000 <= Struct24 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct29 x_10 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_000_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_000_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_000_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_000_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_000(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_000_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_000);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_000);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_000);
        Struct25 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_000 <= (Bit#(2))'(2'h3);
        readLine_000 <= (x_4).victim_line;

        end else begin

            Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_000 <= (Bit#(2))'(2'h3);
                readLine_000 <= (x_5).victim_line;

            end else begin

                Struct25 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_000 <= (Bit#(2))'(2'h3);
                    readLine_000 <= (x_6).victim_line;

                end else begin

                    Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_000 <= (Bit#(2))'(2'h3);
                        readLine_000 <= (x_7).victim_line;

                    end else begin

                        readStage_000 <= (Bit#(2))'(2'h1);
                        readAddr_000 <= x_0;
                        Bit#(8) x_8 = ((x_0)[12:5]);
                        Struct29 x_9 = (Struct29 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_000_0(x_9);
                        let x_11 <- putRq_infoRam_000_1(x_9);
                        let x_12 <- putRq_infoRam_000_2(x_9);
                        let x_13 <- putRq_infoRam_000_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_000_readRs ();
        let x_1 = (readStage_000);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_000 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_000);
        return x_2;
    endmethod

    method Action cache_000_writeRq (Struct24 x_0);
        let x_1 = (readStage_000);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_000);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_000);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct24 x_6 = (Struct24 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_000 <= x_6;
            victims_000 <= update (x_3, (Bit#(2))'(2'h0), Struct25
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct24 x_8 = (Struct24 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_000 <= x_8;
                victims_000 <= update (x_3, (Bit#(2))'(2'h1), Struct25
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct25 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct24 x_10 = (Struct24 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_000 <= x_10;
                    victims_000 <= update (x_3, (Bit#(2))'(2'h2), Struct25
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct25 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct24 x_12 = (Struct24 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_000 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_000 <= x_12;
                        victims_000 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct25 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin
                    writeStage_000 <= (Bit#(3))'(3'h1);
                    writeLine_000 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_000_writeRs ();
        let x_1 = (writeStage_000);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_000 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_000);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_000_hasVictimSlot ();
        let x_1 = (victims_000);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct24) cache_000_getVictim ();
        let x_1 = (victims_000);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct24 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_000_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_000);
        Struct25 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_000 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


        end else begin

            Struct25 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_000 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


            end else begin

                Struct25 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_000 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                end else begin

                    Struct25 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_000 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module66; method Action makeEnq_parentChildren000 (Struct10 x_0);

endinterface


module mkModule66#(function Action enq_fifo00002(Struct2 _),
  function Action enq_fifo0001(Struct2 _),
  function Action enq_fifo0000(Struct2 _)) (Module66);

    // No rules in this module

    method Action makeEnq_parentChildren000 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo0000((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo0001((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo00002(x_3);

            end

        end

    endmethod

endmodule

interface Module67;
    method Action cache_001_readRq (Bit#(64) x_0);
    method ActionValue#(Struct24) cache_001_readRs ();
    method Action cache_001_writeRq (Struct24 x_0);
    method ActionValue#(Struct24) cache_001_writeRs ();
    method ActionValue#(Bool) cache_001_hasVictimSlot ();
    method ActionValue#(Struct24) cache_001_getVictim ();
    method Action cache_001_removeVictim (Bit#(64) x_0);

endinterface


module mkModule67#(function Action putRq_infoRam_001_3(Struct29 _),
  function Action putRq_infoRam_001_2(Struct29 _),
  function Action putRq_infoRam_001_1(Struct29 _),
  function Action putRq_infoRam_001_0(Struct29 _),
  function ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_001(),
  function Action putRq_dataRam_001(Struct28 _),
  function ActionValue#(Struct26) getRs_infoRam_001_3(),
  function ActionValue#(Struct26) getRs_infoRam_001_2(),
  function ActionValue#(Struct26) getRs_infoRam_001_1(),
  function ActionValue#(Struct26) getRs_infoRam_001_0()) (Module67);
    Reg#(Bit#(2)) readStage_001 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_001 <- mkReg(unpack(0));
    Reg#(Struct24) readLine_001 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_001 <- mkReg(unpack(0));
    Reg#(Struct24) writeLine_001 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct25)) victims_001 <- mkReg(unpack(0));
    Reg#(Struct24) victimLine_001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_001 <- mkReg(unpack(0));

    rule read_tagmatch_001;
        let x_0 = (readStage_001);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_001);
        Bit#(51) x_2 = ((x_1)[63:13]);
        Bit#(8) x_3 = ((x_1)[12:5]);
        Vector#(4, Struct26) x_4 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_001_0();
        Vector#(4, Struct26) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_001_1();
        Vector#(4, Struct26) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_001_2();
        Vector#(4, Struct26) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_001_3();
        Vector#(4, Struct26) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct27 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct27 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct27)'(Struct27 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_001 <= Struct24 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        if ((x_13).tm_hit) begin

            readStage_001 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_001(Struct28 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain :
            (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

        end else begin
        readStage_001 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_001;
        let x_0 = (readStage_001);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_001 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_001();
        let x_2 = (readLine_001);
        readLine_001 <= Struct24 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_001);
        when ((x_1).info_hit, noAction);
        writeStage_001 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct29 x_6 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_001_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_001_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_001_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_001_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_001(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_001);
        when (! ((x_1).info_hit), noAction);
        writeStage_001 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Struct29 x_4 = (Struct29 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_001_0(x_4);
        let x_6 <- putRq_infoRam_001_1(x_4);
        let x_7 <- putRq_infoRam_001_2(x_4);
        let x_8 <- putRq_infoRam_001_3(x_4);

    endrule

    rule write_info_miss_rep_rs_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_001 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct26) x_1 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_001_0();
        Vector#(4, Struct26) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_001_1();
        Vector#(4, Struct26) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_001_2();
        Vector#(4, Struct26) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_001_3();
        Vector#(4, Struct26) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_001);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(8) x_13 = ((x_12)[12:5]);
        Struct26 x_14 = ((x_9)[x_10]);
        Bit#(51) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_001 <= x_10;
        victimLine_001 <= Struct24 {addr :
        {(x_15),({(x_13),((Bit#(5))'(5'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        let x_17 <- putRq_dataRam_001(Struct28 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

    endrule

    rule write_victim_rs_001;
        let x_0 = (writeStage_001);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_001);
        writeStage_001 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        let x_5 = (victimWay_001);
        let x_6 = (victims_001);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_001();
        let x_9 = (victimLine_001);
        victims_001 <= update (x_6, x_7, Struct25 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct24 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_001 <= Struct24 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct29 x_10 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_001_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_001_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_001_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_001_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_001(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_001_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_001);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_001);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_001);
        Struct25 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_001 <= (Bit#(2))'(2'h3);
        readLine_001 <= (x_4).victim_line;

        end else begin

            Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_001 <= (Bit#(2))'(2'h3);
                readLine_001 <= (x_5).victim_line;

            end else begin

                Struct25 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_001 <= (Bit#(2))'(2'h3);
                    readLine_001 <= (x_6).victim_line;

                end else begin

                    Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_001 <= (Bit#(2))'(2'h3);
                        readLine_001 <= (x_7).victim_line;

                    end else begin

                        readStage_001 <= (Bit#(2))'(2'h1);
                        readAddr_001 <= x_0;
                        Bit#(8) x_8 = ((x_0)[12:5]);
                        Struct29 x_9 = (Struct29 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_001_0(x_9);
                        let x_11 <- putRq_infoRam_001_1(x_9);
                        let x_12 <- putRq_infoRam_001_2(x_9);
                        let x_13 <- putRq_infoRam_001_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_001_readRs ();
        let x_1 = (readStage_001);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_001 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_001);
        return x_2;
    endmethod

    method Action cache_001_writeRq (Struct24 x_0);
        let x_1 = (readStage_001);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_001);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_001);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct24 x_6 = (Struct24 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_001 <= x_6;
            victims_001 <= update (x_3, (Bit#(2))'(2'h0), Struct25
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct24 x_8 = (Struct24 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_001 <= x_8;
                victims_001 <= update (x_3, (Bit#(2))'(2'h1), Struct25
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct25 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct24 x_10 = (Struct24 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_001 <= x_10;
                    victims_001 <= update (x_3, (Bit#(2))'(2'h2), Struct25
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct25 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct24 x_12 = (Struct24 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_001 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_001 <= x_12;
                        victims_001 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct25 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin
                    writeStage_001 <= (Bit#(3))'(3'h1);
                    writeLine_001 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_001_writeRs ();
        let x_1 = (writeStage_001);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_001 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_001);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_001_hasVictimSlot ();
        let x_1 = (victims_001);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct24) cache_001_getVictim ();
        let x_1 = (victims_001);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct24 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_001_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_001);
        Struct25 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_001 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


        end else begin

            Struct25 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_001 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


            end else begin

                Struct25 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_001 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                end else begin

                    Struct25 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_001 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module68; method Action makeEnq_parentChildren001 (Struct10 x_0);

endinterface


module mkModule68#(function Action enq_fifo00102(Struct2 _),
  function Action enq_fifo0011(Struct2 _),
  function Action enq_fifo0010(Struct2 _)) (Module68);

    // No rules in this module

    method Action makeEnq_parentChildren001 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo0010((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo0011((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo00102(x_3);

            end

        end

    endmethod

endmodule

interface Module69;
    method Action cache_002_readRq (Bit#(64) x_0);
    method ActionValue#(Struct24) cache_002_readRs ();
    method Action cache_002_writeRq (Struct24 x_0);
    method ActionValue#(Struct24) cache_002_writeRs ();
    method ActionValue#(Bool) cache_002_hasVictimSlot ();
    method ActionValue#(Struct24) cache_002_getVictim ();
    method Action cache_002_removeVictim (Bit#(64) x_0);

endinterface


module mkModule69#(function Action putRq_infoRam_002_3(Struct29 _),
  function Action putRq_infoRam_002_2(Struct29 _),
  function Action putRq_infoRam_002_1(Struct29 _),
  function Action putRq_infoRam_002_0(Struct29 _),
  function ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_002(),
  function Action putRq_dataRam_002(Struct28 _),
  function ActionValue#(Struct26) getRs_infoRam_002_3(),
  function ActionValue#(Struct26) getRs_infoRam_002_2(),
  function ActionValue#(Struct26) getRs_infoRam_002_1(),
  function ActionValue#(Struct26) getRs_infoRam_002_0()) (Module69);
    Reg#(Bit#(2)) readStage_002 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_002 <- mkReg(unpack(0));
    Reg#(Struct24) readLine_002 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_002 <- mkReg(unpack(0));
    Reg#(Struct24) writeLine_002 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct25)) victims_002 <- mkReg(unpack(0));
    Reg#(Struct24) victimLine_002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_002 <- mkReg(unpack(0));

    rule read_tagmatch_002;
        let x_0 = (readStage_002);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_002);
        Bit#(51) x_2 = ((x_1)[63:13]);
        Bit#(8) x_3 = ((x_1)[12:5]);
        Vector#(4, Struct26) x_4 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_002_0();
        Vector#(4, Struct26) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_002_1();
        Vector#(4, Struct26) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_002_2();
        Vector#(4, Struct26) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_002_3();
        Vector#(4, Struct26) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct27 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct27 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct27)'(Struct27 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_002 <= Struct24 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        if ((x_13).tm_hit) begin

            readStage_002 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_002(Struct28 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain :
            (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

        end else begin
        readStage_002 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_002;
        let x_0 = (readStage_002);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_002 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_002();
        let x_2 = (readLine_002);
        readLine_002 <= Struct24 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_002;
        let x_0 = (writeStage_002);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_002);
        when ((x_1).info_hit, noAction);
        writeStage_002 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct29 x_6 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_002_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_002_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_002_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_002_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_002(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_002;
        let x_0 = (writeStage_002);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_002);
        when (! ((x_1).info_hit), noAction);
        writeStage_002 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Struct29 x_4 = (Struct29 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_002_0(x_4);
        let x_6 <- putRq_infoRam_002_1(x_4);
        let x_7 <- putRq_infoRam_002_2(x_4);
        let x_8 <- putRq_infoRam_002_3(x_4);

    endrule

    rule write_info_miss_rep_rs_002;
        let x_0 = (writeStage_002);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_002 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct26) x_1 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_002_0();
        Vector#(4, Struct26) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_002_1();
        Vector#(4, Struct26) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_002_2();
        Vector#(4, Struct26) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_002_3();
        Vector#(4, Struct26) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_002);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(8) x_13 = ((x_12)[12:5]);
        Struct26 x_14 = ((x_9)[x_10]);
        Bit#(51) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_002 <= x_10;
        victimLine_002 <= Struct24 {addr :
        {(x_15),({(x_13),((Bit#(5))'(5'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        let x_17 <- putRq_dataRam_002(Struct28 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

    endrule

    rule write_victim_rs_002;
        let x_0 = (writeStage_002);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_002);
        writeStage_002 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        let x_5 = (victimWay_002);
        let x_6 = (victims_002);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_002();
        let x_9 = (victimLine_002);
        victims_002 <= update (x_6, x_7, Struct25 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct24 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_002 <= Struct24 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct29 x_10 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_002_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_002_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_002_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_002_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_002(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_002_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_002);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_002);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_002);
        Struct25 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_002 <= (Bit#(2))'(2'h3);
        readLine_002 <= (x_4).victim_line;

        end else begin

            Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_002 <= (Bit#(2))'(2'h3);
                readLine_002 <= (x_5).victim_line;

            end else begin

                Struct25 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_002 <= (Bit#(2))'(2'h3);
                    readLine_002 <= (x_6).victim_line;

                end else begin

                    Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_002 <= (Bit#(2))'(2'h3);
                        readLine_002 <= (x_7).victim_line;

                    end else begin

                        readStage_002 <= (Bit#(2))'(2'h1);
                        readAddr_002 <= x_0;
                        Bit#(8) x_8 = ((x_0)[12:5]);
                        Struct29 x_9 = (Struct29 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_002_0(x_9);
                        let x_11 <- putRq_infoRam_002_1(x_9);
                        let x_12 <- putRq_infoRam_002_2(x_9);
                        let x_13 <- putRq_infoRam_002_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_002_readRs ();
        let x_1 = (readStage_002);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_002 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_002);
        return x_2;
    endmethod

    method Action cache_002_writeRq (Struct24 x_0);
        let x_1 = (readStage_002);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_002);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_002);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct24 x_6 = (Struct24 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_002 <= x_6;
            victims_002 <= update (x_3, (Bit#(2))'(2'h0), Struct25
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct24 x_8 = (Struct24 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_002 <= x_8;
                victims_002 <= update (x_3, (Bit#(2))'(2'h1), Struct25
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct25 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct24 x_10 = (Struct24 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_002 <= x_10;
                    victims_002 <= update (x_3, (Bit#(2))'(2'h2), Struct25
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct25 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct24 x_12 = (Struct24 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_002 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_002 <= x_12;
                        victims_002 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct25 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin
                    writeStage_002 <= (Bit#(3))'(3'h1);
                    writeLine_002 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_002_writeRs ();
        let x_1 = (writeStage_002);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_002 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_002);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_002_hasVictimSlot ();
        let x_1 = (victims_002);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct24) cache_002_getVictim ();
        let x_1 = (victims_002);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct24 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_002_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_002);
        Struct25 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_002 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


        end else begin

            Struct25 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_002 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


            end else begin

                Struct25 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_002 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                end else begin

                    Struct25 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_002 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module70; method Action makeEnq_parentChildren002 (Struct10 x_0);

endinterface


module mkModule70#(function Action enq_fifo00202(Struct2 _),
  function Action enq_fifo0021(Struct2 _),
  function Action enq_fifo0020(Struct2 _)) (Module70);

    // No rules in this module

    method Action makeEnq_parentChildren002 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo0020((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo0021((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo00202(x_3);

            end

        end

    endmethod

endmodule

interface Module71;
    method Action cache_003_readRq (Bit#(64) x_0);
    method ActionValue#(Struct24) cache_003_readRs ();
    method Action cache_003_writeRq (Struct24 x_0);
    method ActionValue#(Struct24) cache_003_writeRs ();
    method ActionValue#(Bool) cache_003_hasVictimSlot ();
    method ActionValue#(Struct24) cache_003_getVictim ();
    method Action cache_003_removeVictim (Bit#(64) x_0);

endinterface


module mkModule71#(function Action putRq_infoRam_003_3(Struct29 _),
  function Action putRq_infoRam_003_2(Struct29 _),
  function Action putRq_infoRam_003_1(Struct29 _),
  function Action putRq_infoRam_003_0(Struct29 _),
  function ActionValue#(Vector#(4, Bit#(64))) getRs_dataRam_003(),
  function Action putRq_dataRam_003(Struct28 _),
  function ActionValue#(Struct26) getRs_infoRam_003_3(),
  function ActionValue#(Struct26) getRs_infoRam_003_2(),
  function ActionValue#(Struct26) getRs_infoRam_003_1(),
  function ActionValue#(Struct26) getRs_infoRam_003_0()) (Module71);
    Reg#(Bit#(2)) readStage_003 <- mkReg(unpack(0));
    Reg#(Bit#(64)) readAddr_003 <- mkReg(unpack(0));
    Reg#(Struct24) readLine_003 <- mkReg(unpack(0));
    Reg#(Bit#(3)) writeStage_003 <- mkReg(unpack(0));
    Reg#(Struct24) writeLine_003 <- mkReg(unpack(0));
    Reg#(Vector#(4, Struct25)) victims_003 <- mkReg(unpack(0));
    Reg#(Struct24) victimLine_003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) victimWay_003 <- mkReg(unpack(0));

    rule read_tagmatch_003;
        let x_0 = (readStage_003);
        when ((x_0) == ((Bit#(2))'(2'h1)), noAction);
        let x_1 = (readAddr_003);
        Bit#(51) x_2 = ((x_1)[63:13]);
        Bit#(8) x_3 = ((x_1)[12:5]);
        Vector#(4, Struct26) x_4 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_5 <- getRs_infoRam_003_0();
        Vector#(4, Struct26) x_6 = (update (x_4, (Bit#(2))'(2'h0), x_5));
        let x_7 <- getRs_infoRam_003_1();
        Vector#(4, Struct26) x_8 = (update (x_6, (Bit#(2))'(2'h1), x_7));
        let x_9 <- getRs_infoRam_003_2();
        Vector#(4, Struct26) x_10 = (update (x_8, (Bit#(2))'(2'h2), x_9));
        let x_11 <- getRs_infoRam_003_3();
        Vector#(4, Struct26) x_12 = (update (x_10, (Bit#(2))'(2'h3), x_11));

        Struct27 x_13 = (((((x_12)[(Bit#(2))'(2'h0)]).tag) == (x_2) ?
        (Struct27 {tm_hit : (Bool)'(True), tm_way : (Bit#(2))'(2'h0),
        tm_value : ((x_12)[(Bit#(2))'(2'h0)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h1)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h1), tm_value :
        ((x_12)[(Bit#(2))'(2'h1)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h2)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h2), tm_value :
        ((x_12)[(Bit#(2))'(2'h2)]).value}) :
        (((((x_12)[(Bit#(2))'(2'h3)]).tag) == (x_2) ? (Struct27 {tm_hit :
        (Bool)'(True), tm_way : (Bit#(2))'(2'h3), tm_value :
        ((x_12)[(Bit#(2))'(2'h3)]).value}) :
        ((Struct27)'(Struct27 {tm_hit: False, tm_way: 2'h0, tm_value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}))))))))));

        readLine_003 <= Struct24 {addr : x_1, info_hit : (x_13).tm_hit,
        info_way : (x_13).tm_way, info_write : (Bool)'(False), info :
        (x_13).tm_value, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        if ((x_13).tm_hit) begin

            readStage_003 <= (Bit#(2))'(2'h2);
            let x_14 <- putRq_dataRam_003(Struct28 {write : (Bool)'(False),
            addr : {(x_3),((x_13).tm_way)}, datain :
            (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

        end else begin
        readStage_003 <= (Bit#(2))'(2'h3);

        end

    endrule

    rule read_data_003;
        let x_0 = (readStage_003);
        when ((x_0) == ((Bit#(2))'(2'h2)), noAction);
        readStage_003 <= (Bit#(2))'(2'h3);
        let x_1 <- getRs_dataRam_003();
        let x_2 = (readLine_003);
        readLine_003 <= Struct24 {addr : (x_2).addr, info_hit :
        (x_2).info_hit, info_way : (x_2).info_way, info_write :
        (x_2).info_write, info : (x_2).info, value_write : (Bool)'(False),
        value : x_1};

    endrule

    rule write_info_hit_003;
        let x_0 = (writeStage_003);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_003);
        when ((x_1).info_hit, noAction);
        writeStage_003 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        Bit#(2) x_5 = ((x_1).info_way);
        if ((x_1).info_write) begin

            Struct29 x_6 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_7 <- putRq_infoRam_003_0(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_9 <- putRq_infoRam_003_1(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_11 <- putRq_infoRam_003_2(x_6);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_13 <- putRq_infoRam_003_3(x_6);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_16 <- putRq_dataRam_003(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule

    rule write_info_miss_rep_rq_003;
        let x_0 = (writeStage_003);
        when ((x_0) == ((Bit#(3))'(3'h1)), noAction);
        let x_1 = (writeLine_003);
        when (! ((x_1).info_hit), noAction);
        writeStage_003 <= (Bit#(3))'(3'h2);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(8) x_3 = ((x_2)[12:5]);
        Struct29 x_4 = (Struct29 {write : (Bool)'(False), addr : x_3, datain
        :
        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

        let x_5 <- putRq_infoRam_003_0(x_4);
        let x_6 <- putRq_infoRam_003_1(x_4);
        let x_7 <- putRq_infoRam_003_2(x_4);
        let x_8 <- putRq_infoRam_003_3(x_4);

    endrule

    rule write_info_miss_rep_rs_003;
        let x_0 = (writeStage_003);
        when ((x_0) == ((Bit#(3))'(3'h2)), noAction);
        writeStage_003 <= (Bit#(3))'(3'h3);
        Vector#(4, Struct26) x_1 =
        ((Vector#(4, Struct26))'(vec(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}}, Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})));

        let x_2 <- getRs_infoRam_003_0();
        Vector#(4, Struct26) x_3 = (update (x_1, (Bit#(2))'(2'h0), x_2));
        let x_4 <- getRs_infoRam_003_1();
        Vector#(4, Struct26) x_5 = (update (x_3, (Bit#(2))'(2'h1), x_4));
        let x_6 <- getRs_infoRam_003_2();
        Vector#(4, Struct26) x_7 = (update (x_5, (Bit#(2))'(2'h2), x_6));
        let x_8 <- getRs_infoRam_003_3();
        Vector#(4, Struct26) x_9 = (update (x_7, (Bit#(2))'(2'h3), x_8));

        Bit#(2) x_10 = ((((((x_9)[(Bit#(2))'(2'h0)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h0)) :
        ((((((x_9)[(Bit#(2))'(2'h1)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h1)) :
        ((((((x_9)[(Bit#(2))'(2'h2)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h2)) :
        ((((((x_9)[(Bit#(2))'(2'h3)]).value).mesi_dir_st) ==
        ((Bit#(3))'(3'h1)) ? ((Bit#(2))'(2'h3)) : ((Bit#(2))'(2'h0))))))))));

        let x_11 = (writeLine_003);
        Bit#(64) x_12 = ((x_11).addr);
        Bit#(8) x_13 = ((x_12)[12:5]);
        Struct26 x_14 = ((x_9)[x_10]);
        Bit#(51) x_15 = ((x_14).tag);
        Struct4 x_16 = ((x_14).value);
        victimWay_003 <= x_10;
        victimLine_003 <= Struct24 {addr :
        {(x_15),({(x_13),((Bit#(5))'(5'h0))})}, info_hit : (Bool)'(False),
        info_way : (Bit#(2))'(2'h0), info_write : (Bool)'(False), info :
        x_16, value_write : (Bool)'(False), value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))};
        let x_17 <- putRq_dataRam_003(Struct28 {write : (Bool)'(False), addr
        : {(x_13),(x_10)}, datain :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});

    endrule

    rule write_victim_rs_003;
        let x_0 = (writeStage_003);
        when ((x_0) == ((Bit#(3))'(3'h3)), noAction);
        let x_1 = (writeLine_003);
        writeStage_003 <= (Bit#(3))'(3'h7);
        Bit#(64) x_2 = ((x_1).addr);
        Bit#(51) x_3 = ((x_2)[63:13]);
        Bit#(8) x_4 = ((x_2)[12:5]);
        let x_5 = (victimWay_003);
        let x_6 = (victims_003);
        when ((! (((x_6)[(Bit#(2))'(2'h3)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h2)]).victim_valid)) || ((!
        (((x_6)[(Bit#(2))'(2'h1)]).victim_valid)) || (!
        (((x_6)[(Bit#(2))'(2'h0)]).victim_valid)))), noAction);
        Bit#(2) x_7 = ((((x_6)[(Bit#(2))'(2'h3)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h2)]).victim_valid ?
        ((((x_6)[(Bit#(2))'(2'h1)]).victim_valid ? ((Bit#(2))'(2'h0)) :
        ((Bit#(2))'(2'h1)))) : ((Bit#(2))'(2'h2)))) : ((Bit#(2))'(2'h3))));

        let x_8 <- getRs_dataRam_003();
        let x_9 = (victimLine_003);
        victims_003 <= update (x_6, x_7, Struct25 {victim_valid :
        (Bool)'(True), victim_idx : x_7, victim_line : Struct24 {addr :
        (x_9).addr, info_hit : (x_9).info_hit, info_way : (x_9).info_way,
        info_write : (x_9).info_write, info : (x_9).info, value_write :
        (Bool)'(False), value : x_8}});
        writeLine_003 <= Struct24 {addr : x_2, info_hit : (Bool)'(True),
        info_way : x_5, info_write : (Bool)'(False), info : (x_1).info,
        value_write : (Bool)'(False), value : (x_1).value};
        if ((x_1).info_write) begin

            Struct29 x_10 = (Struct29 {write : (Bool)'(True), addr : x_4,
            datain : Struct26 {tag : x_3, value : (x_1).info}});
            if ((x_5) == ((Bit#(2))'(2'h0))) begin
            let x_11 <- putRq_infoRam_003_0(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h1))) begin
            let x_13 <- putRq_infoRam_003_1(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h2))) begin
            let x_15 <- putRq_infoRam_003_2(x_10);

            end else begin

            end
            if ((x_5) == ((Bit#(2))'(2'h3))) begin
            let x_17 <- putRq_infoRam_003_3(x_10);

            end else begin

            end

        end else begin

        end
        if ((x_1).value_write) begin

            let x_20 <- putRq_dataRam_003(Struct28 {write : (Bool)'(True),
            addr : {(x_4),(x_5)}, datain : (x_1).value});

        end else begin

        end

    endrule


    method Action cache_003_readRq (Bit#(64) x_0);
        let x_1 = (writeStage_003);
        when ((x_1) == ((Bit#(3))'(3'h0)), noAction);
        let x_2 = (readStage_003);
        when ((x_2) == ((Bit#(2))'(2'h0)), noAction);
        let x_3 = (victims_003);
        Struct25 x_4 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_4).victim_valid) && ((((x_4).victim_line).addr) == (x_0)))
        begin
        readStage_003 <= (Bit#(2))'(2'h3);
        readLine_003 <= (x_4).victim_line;

        end else begin

            Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
            (x_0))) begin

                readStage_003 <= (Bit#(2))'(2'h3);
                readLine_003 <= (x_5).victim_line;

            end else begin

                Struct25 x_6 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_6).victim_valid) && ((((x_6).victim_line).addr) ==
                (x_0))) begin

                    readStage_003 <= (Bit#(2))'(2'h3);
                    readLine_003 <= (x_6).victim_line;

                end else begin

                    Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_7).victim_valid) && ((((x_7).victim_line).addr)
                    == (x_0))) begin

                        readStage_003 <= (Bit#(2))'(2'h3);
                        readLine_003 <= (x_7).victim_line;

                    end else begin

                        readStage_003 <= (Bit#(2))'(2'h1);
                        readAddr_003 <= x_0;
                        Bit#(8) x_8 = ((x_0)[12:5]);
                        Struct29 x_9 = (Struct29 {write : (Bool)'(False),
                        addr : x_8, datain :
                        (Struct26)'(Struct26 {tag: 51'h0, value: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}})});

                        let x_10 <- putRq_infoRam_003_0(x_9);
                        let x_11 <- putRq_infoRam_003_1(x_9);
                        let x_12 <- putRq_infoRam_003_2(x_9);
                        let x_13 <- putRq_infoRam_003_3(x_9);

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_003_readRs ();
        let x_1 = (readStage_003);
        when ((x_1) == ((Bit#(2))'(2'h3)), noAction);
        readStage_003 <= (Bit#(2))'(2'h0);
        let x_2 = (readLine_003);
        return x_2;
    endmethod

    method Action cache_003_writeRq (Struct24 x_0);
        let x_1 = (readStage_003);
        when ((x_1) == ((Bit#(2))'(2'h0)), noAction);
        let x_2 = (writeStage_003);
        when ((x_2) == ((Bit#(3))'(3'h0)), noAction);
        let x_3 = (victims_003);
        Bool x_4 = ((((x_0).info).mesi_dir_st) == ((Bit#(3))'(3'h1)));

        Struct25 x_5 = ((x_3)[(Bit#(2))'(2'h0)]);
        if (((x_5).victim_valid) && ((((x_5).victim_line).addr) ==
        ((x_0).addr))) begin

            Struct24 x_6 = (Struct24 {addr : (x_0).addr, info_hit :
            (Bool)'(False), info_way : (x_0).info_way, info_write :
            (x_0).info_write, info : (x_0).info, value_write :
            (x_0).value_write, value : (x_0).value});
            writeStage_003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
            ((Bit#(3))'(3'h1)));
            writeLine_003 <= x_6;
            victims_003 <= update (x_3, (Bit#(2))'(2'h0), Struct25
            {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h0), victim_line :
            x_6});

        end else begin

            Struct25 x_7 = ((x_3)[(Bit#(2))'(2'h1)]);
            if (((x_7).victim_valid) && ((((x_7).victim_line).addr) ==
            ((x_0).addr))) begin

                Struct24 x_8 = (Struct24 {addr : (x_0).addr, info_hit :
                (Bool)'(False), info_way : (x_0).info_way, info_write :
                (x_0).info_write, info : (x_0).info, value_write :
                (x_0).value_write, value : (x_0).value});
                writeStage_003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                ((Bit#(3))'(3'h1)));
                writeLine_003 <= x_8;
                victims_003 <= update (x_3, (Bit#(2))'(2'h1), Struct25
                {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h1),
                victim_line : x_8});

            end else begin

                Struct25 x_9 = ((x_3)[(Bit#(2))'(2'h2)]);
                if (((x_9).victim_valid) && ((((x_9).victim_line).addr) ==
                ((x_0).addr))) begin

                    Struct24 x_10 = (Struct24 {addr : (x_0).addr, info_hit :
                    (Bool)'(False), info_way : (x_0).info_way, info_write :
                    (x_0).info_write, info : (x_0).info, value_write :
                    (x_0).value_write, value : (x_0).value});
                    writeStage_003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                    ((Bit#(3))'(3'h1)));
                    writeLine_003 <= x_10;
                    victims_003 <= update (x_3, (Bit#(2))'(2'h2), Struct25
                    {victim_valid : x_4, victim_idx : (Bit#(2))'(2'h2),
                    victim_line : x_10});

                end else begin

                    Struct25 x_11 = ((x_3)[(Bit#(2))'(2'h3)]);
                    if (((x_11).victim_valid) && ((((x_11).victim_line).addr)
                    == ((x_0).addr))) begin

                        Struct24 x_12 = (Struct24 {addr : (x_0).addr,
                        info_hit : (Bool)'(False), info_way : (x_0).info_way,
                        info_write : (x_0).info_write, info : (x_0).info,
                        value_write : (x_0).value_write, value :
                        (x_0).value});
                        writeStage_003 <= (x_4 ? ((Bit#(3))'(3'h7)) :
                        ((Bit#(3))'(3'h1)));
                        writeLine_003 <= x_12;
                        victims_003 <= update (x_3, (Bit#(2))'(2'h3),
                        Struct25 {victim_valid : x_4, victim_idx :
                        (Bit#(2))'(2'h3), victim_line : x_12});

                    end else begin
                    writeStage_003 <= (Bit#(3))'(3'h1);
                    writeLine_003 <= x_0;

                    end

                end

            end

        end

    endmethod

    method ActionValue#(Struct24) cache_003_writeRs ();
        let x_1 = (writeStage_003);
        when ((x_1) == ((Bit#(3))'(3'h7)), noAction);
        writeStage_003 <= (Bit#(3))'(3'h0);
        let x_2 = (writeLine_003);
        return x_2;
    endmethod

    method ActionValue#(Bool) cache_003_hasVictimSlot ();
        let x_1 = (victims_003);
        Bool x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))));
        return x_2;
    endmethod

    method ActionValue#(Struct24) cache_003_getVictim ();
        let x_1 = (victims_003);
        when ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid) ||
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid) ||
        (((x_1)[(Bit#(2))'(2'h0)]).victim_valid))), noAction);
        Struct24 x_2 = ((((x_1)[(Bit#(2))'(2'h3)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h3)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h2)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h2)]).victim_line) :
        ((((x_1)[(Bit#(2))'(2'h1)]).victim_valid ?
        (((x_1)[(Bit#(2))'(2'h1)]).victim_line) :
        (((x_1)[(Bit#(2))'(2'h0)]).victim_line)))))));
        return x_2;
    endmethod

    method Action cache_003_removeVictim (Bit#(64) x_0);
        let x_1 = (victims_003);
        Struct25 x_2 = ((x_1)[(Bit#(2))'(2'h0)]);
        if (((x_2).victim_valid) && ((((x_2).victim_line).addr) == (x_0)))
        begin

            victims_003 <= update (x_1, (Bit#(2))'(2'h0),
            (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


        end else begin

            Struct25 x_3 = ((x_1)[(Bit#(2))'(2'h1)]);
            if (((x_3).victim_valid) && ((((x_3).victim_line).addr) ==
            (x_0))) begin

                victims_003 <= update (x_1, (Bit#(2))'(2'h1),
                (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


            end else begin

                Struct25 x_4 = ((x_1)[(Bit#(2))'(2'h2)]);
                if (((x_4).victim_valid) && ((((x_4).victim_line).addr) ==
                (x_0))) begin

                    victims_003 <= update (x_1, (Bit#(2))'(2'h2),
                    (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                end else begin

                    Struct25 x_5 = ((x_1)[(Bit#(2))'(2'h3)]);
                    if (((x_5).victim_valid) && ((((x_5).victim_line).addr)
                    == (x_0))) begin

                        victims_003 <= update (x_1, (Bit#(2))'(2'h3),
                        (Struct25)'(Struct25 {victim_valid: False, victim_idx: 2'h0, victim_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}}));


                    end else begin

                    end

                end

            end

        end

    endmethod

endmodule

interface Module72; method Action makeEnq_parentChildren003 (Struct10 x_0);

endinterface


module mkModule72#(function Action enq_fifo00302(Struct2 _),
  function Action enq_fifo0031(Struct2 _),
  function Action enq_fifo0030(Struct2 _)) (Module72);

    // No rules in this module

    method Action makeEnq_parentChildren003 (Struct10 x_0);
        if (((x_0).enq_type) == ((Bit#(2))'(2'h0))) begin
        let x_1 <- enq_fifo0030((x_0).enq_msg);

        end else begin

            if (((x_0).enq_type) == ((Bit#(2))'(2'h1))) begin
            let x_2 <- enq_fifo0031((x_0).enq_msg);

            end else begin
            Struct2 x_3 = ((x_0).enq_msg);
            let x_4 <- enq_fifo00302(x_3);

            end

        end

    endmethod

endmodule

interface Module73;
endinterface


module mkModule73#(function ActionValue#(Struct3) cache_00_writeRs(),
  function Action cache_00_removeVictim(Bit#(64) _),
  function ActionValue#(Struct3) cache_00_getVictim(),
  function Action transferUpDown00(Struct17 _),
  function Action releaseDL00(Bit#(64) _),
  function Action releaseUL00(Bit#(64) _),
  function ActionValue#(Struct15) upLockGet00(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0031(),
  function ActionValue#(Struct2) deq_fifo0021(),
  function ActionValue#(Struct2) deq_fifo0011(),
  function Action addRs00(Struct14 _),
  function ActionValue#(Struct6) downLockGet00(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0001(),
  function Action broadcast_parentChildren00(Struct13 _),
  function Action registerDL00(Struct12 _),
  function Action registerUL00(Struct11 _),
  function ActionValue#(Bool) cache_00_hasVictimSlot(),
  function Action makeEnq_parentChildren00(Struct10 _),
  function Action cache_00_writeRq(Struct3 _),
  function ActionValue#(Bool) downLockable00(Bit#(64) _),
  function ActionValue#(Bool) upLockable00(Bit#(64) _),
  function ActionValue#(Struct3) cache_00_readRs(),
  function ActionValue#(Struct2) deq_fifo0030(),
  function ActionValue#(Struct2) deq_fifo0020(),
  function ActionValue#(Struct2) deq_fifo0010(),
  function ActionValue#(Struct2) deq_fifo0000(),
  function ActionValue#(Struct6) downLockRssFull00(),
  function Action cache_00_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo002()) (Module73);
    Reg#(Bit#(1)) rr00 <- mkReg(unpack(0));
    Reg#(Struct1) prl00 <- mkReg(unpack(0));
    Reg#(Struct1) crqrl00 <- mkReg(unpack(0));
    Reg#(Struct1) crsrl00 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc00 <- mkReg(unpack(0));
    Reg#(Struct5) wl00 <- mkReg(unpack(0));

    rule rr_00;let x_0 = (rr00);
               rr00 <= (x_0) + ((Bit#(1))'(1'h1));

    endrule

    rule rule_00_1230;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo002();
        prl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc00 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_1232;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull00();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc00 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_00_readRq((x_4).addr);

    endrule

    rule rule_00_12310000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo0000();
        crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc00 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_12310010;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo0010();
        crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h1), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc00 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_12310020;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo0020();
        crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h2), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc00 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_12310030;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo0030();
        crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h3), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc00 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_00_readRq((x_3).addr);

    endrule

    rule rule_00_456;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        let x_3 <- cache_00_readRs();
        let x_4 = (rlc00);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl00 <= Struct1 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl00 <= Struct1 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl00 <= Struct1 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_00_000000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_001000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_01000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_03000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_10000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 = (wl00);
        when (! ((x_23).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_14000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h8)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_15000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))), r_dl_rsbTo : (Bit#(4))'(4'h8)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_25000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_2600000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_2601000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_261000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_27000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_28000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_290000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_291000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_210000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h0))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h0)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_211000;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h0))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h0)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_00_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_040000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0001();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_070000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0001();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1600000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0001();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1601000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0001();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11000000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0001();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11001000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0001();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11002000;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0001();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h4))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_000001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_001001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_01001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_03001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_10001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h1), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 = (wl00);
        when (! ((x_23).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h9))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_14001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h9)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_15001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))), r_dl_rsbTo : (Bit#(4))'(4'h9)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_25001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_2600001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_2601001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_261001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_27001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_28001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_290001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_291001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_210001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h1))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h1)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_211001;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h1)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h1))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h1)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_00_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'h9))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h9))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h9))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_040001;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0011();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_070001;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0011();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1600001;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0011();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1601001;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0011();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11000001;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0011();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11001001;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0011();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11002001;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0011();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h5))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_000002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_001002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_01002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_03002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_10002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h2), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 = (wl00);
        when (! ((x_23).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'ha))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_14002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'ha)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_15002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))), r_dl_rsbTo : (Bit#(4))'(4'ha)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_25002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_2600002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_2601002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_261002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_27002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_28002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_290002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_291002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_210002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h2))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h2)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_211002;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h2)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h2))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h2)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_00_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'ha))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'ha))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'ha))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_040002;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0021();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_070002;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0021();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1600002;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0021();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1601002;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0021();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11000002;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0021();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11001002;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0021();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11002002;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0021();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h6))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_000003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! (((Bit#(3))'(3'h2)) < ((x_10).dir_st))) && ((x_9) ==
        ((Bit#(3))'(3'h2))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) : (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ?
        (((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) :
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))}).dir_excl)))},
        value_write : (x_5).value_write, value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h3), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_001003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h4), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_01003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h1)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_03003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h2)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_10003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) || (((x_9) ==
        ((Bit#(3))'(3'h2))) && (((x_8) == ((Bool)'(True))) &&
        ((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) ==
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (Bit#(2))'(2'h3), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hb), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren00(x_21);
        let x_23 = (wl00);
        when (! ((x_23).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_8) == ((Bool)'(False))) && ((! (((Bit#(3))'(3'h2)) <
        (x_9))) && (! (((Bit#(3))'(3'h2)) < ((x_10).dir_st)))), noAction);

        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_00_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(True), r_ul_msg
        : x_15, r_ul_rsbTo : ((Bit#(4))'(4'hb))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren00(x_18);
        let x_20 = (wl00);
        when (! ((x_20).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_14003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1))
        < (x_9))) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (!
        (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'hb)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_15003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'ha)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))) == ((Bit#(4))'(4'h0)))) && (((x_8) ==
        ((Bool)'(True))) && ((! (((Bit#(3))'(3'h2)) < (x_9))) &&
        (((x_10).dir_st) == ((Bit#(3))'(3'h2))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))), r_dl_rsbTo : (Bit#(4))'(4'hb)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_25003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_2600003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_2601003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_261003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_27003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h14)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h3)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_28003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl)
        == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h1)), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_290003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(False))) && (((((((x_10).dir_st) ==
        ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers))
        ? ((Bit#(3))'(3'h2)) : ((Bit#(3))'(3'h1)))))))) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_291003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((Bit#(3))'(3'h1)) < ((((((x_10).dir_sharers)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((x_10).dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((((((((x_10).dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        (((((((((x_10).dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(3))'(3'h1)) : ((Bit#(3))'(3'h0)))) +
        ((Bit#(3))'(3'h0))))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl,
        dir_sharers : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3))))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_210003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && (((x_9) == ((Bit#(3))'(3'h2))) &&
        (((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ?
        ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) == ((Bit#(3))'(3'h2))) &&
        ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1)) << ((Bit#(2))'(2'h3))))
        == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2)) :
        ((Bit#(3))'(3'h1)))))))) == ((Bit#(3))'(3'h2))) &&
        (((x_10).dir_sharers) == (((Bit#(4))'(4'h1)) <<
        ((Bit#(2))'(2'h3)))))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        let x_19 <- cache_00_writeRq(x_18);
        Struct10 x_20 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_21 <- makeEnq_parentChildren00(x_20);
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_211003;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h3)), noAction);
        Struct3 x_4 = ((x_2).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h15)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable00((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (! ((((((x_10).dir_st) == ((Bit#(3))'(3'h4))) &&
        (((x_10).dir_excl) == ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h4)) :
        (((((x_10).dir_st) == ((Bit#(3))'(3'h3))) && (((x_10).dir_excl) ==
        ((Bit#(2))'(2'h3))) ? ((Bit#(3))'(3'h3)) : (((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && ((((x_10).dir_sharers) | (((Bit#(4))'(4'h1))
        << ((Bit#(2))'(2'h3)))) == ((x_10).dir_sharers)) ? ((Bit#(3))'(3'h2))
        : ((Bit#(3))'(3'h1)))))))) < ((Bit#(3))'(3'h3))), noAction);
        crqrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_19).value_write,
        value : (x_19).value});
        let x_21 <- cache_00_writeRq(x_20);
        Struct10 x_22 = (Struct10 {enq_type : ((((Bit#(4))'(4'hb))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'hb))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'hb))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h16), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_040003;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0031();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_070003;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0031();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'h6)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1600003;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0031();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_1601003;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0031();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11000003;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0031();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11001003;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0031();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hf)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11002003;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        Struct3 x_3 =
        ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}));

        Vector#(4, Bit#(64)) x_4 = ((x_3).value);
        Struct4 x_5 = ((x_3).info);
        Bool x_6 = ((x_5).mesi_owned);
        Bit#(3) x_7 = ((x_5).mesi_status);
        Struct8 x_8 = (Struct8 {dir_st : (x_5).mesi_dir_st, dir_excl :
        ((((x_5).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_5).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_5).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_5).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_5).mesi_dir_sharers});
        let x_9 <- deq_fifo0031();
        Struct9 x_10 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_11 <- downLockGet00((x_9).addr);
        when ((x_11).valid, noAction);
        Struct7 x_12 = ((x_11).data);
        when (((x_9).id) == ((Bit#(6))'(6'hd)), noAction);
        when ((x_12).dl_valid, noAction);
        when ((x_12).dl_rsb, noAction);
        when ((((x_12).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_12).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when ((x_9).type_, noAction);
        when ((Bool)'(True), noAction);
        Struct2 x_13 = (x_9);
        let x_14 <- addRs00(Struct14 {r_dl_addr : (x_9).addr, r_dl_midx :
        ((Bit#(4))'(4'h7))[1:0], r_dl_msg : x_13});
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_020;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_19 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st :
        (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (x_10).dir_excl, dir_sharers :
        (((x_10).dir_st) == ((Bit#(3))'(3'h2)) ? (((x_10).dir_sharers) |
        (((Bit#(4))'(4'h1)) << ((x_18)[1:0]))) : (((Bit#(4))'(4'h1)) <<
        ((x_18)[1:0])))}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct3 x_22 = (Struct3 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_00_writeRq(x_22);
        let x_24 <- releaseUL00((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren00(x_25);
        let x_27 = (wl00);
        when (! ((x_27).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_021;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_19 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h3), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        Struct3 x_22 = (Struct3 {addr : (x_21).addr, info_hit :
        (x_21).info_hit, info_way : (x_21).info_way, info_write :
        (x_21).info_write, info : (x_21).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_23 <- cache_00_writeRq(x_22);
        let x_24 <- releaseUL00((x_11).addr);
        Struct10 x_25 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h4),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_26 <- makeEnq_parentChildren00(x_25);
        let x_27 = (wl00);
        when (! ((x_27).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_041;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h2)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct3 x_18 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_st,
        mesi_dir_sharers : (((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl :
        (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) |
        (((Bit#(4))'(4'h1)) << (((x_15).cidx)[1:0]))}).dir_sharers) :
        (((Bit#(4))'(4'h1)) << ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl
        : (Bit#(2))'(2'h0), dir_sharers : (((Bit#(4))'(4'h0)) |
        (((Bit#(4))'(4'h1)) << ((x_17)[1:0]))) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_00_writeRq(x_21);
        let x_23 <- releaseDL00((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h3),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 = (wl00);
        when (! ((x_26).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_05;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h2)))) && (! (((Bit#(3))'(3'h2)) <
        ((x_10).dir_st))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct3 x_16 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_17 = (Struct3 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_06;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((Bit#(3))'(3'h1)) < (x_9))) && ((!
        (((x_10).dir_st) < ((Bit#(3))'(3'h3)))) && (! (((Bit#(3))'(3'h4)) <
        ((x_10).dir_st))))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'h5), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_071;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'h5)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct16 x_15 = (Struct16 {cidx :
        {((Bit#(2))'(2'h1)),(((((x_14).dl_rss_from)[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))))}, msg :
        ((x_14).dl_rss)[((((x_14).dl_rss_from)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_14).dl_rss_from)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_14).dl_rss_from)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_14).dl_rss_from)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0)))))))))))))]});
        Struct2 x_16 = ((x_14).dl_msg);
        Bit#(4) x_17 = ((x_14).dl_rsbTo);
        Struct3 x_18 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st
        : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8
        {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_sharers) : (((Bit#(4))'(4'h1)) <<
        ((Struct8 {dir_st : (Bit#(3))'(3'h2), dir_excl : (Bit#(2))'(2'h0),
        dir_sharers : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (((x_15).cidx)[1:0]))}).dir_excl)))}, value_write :
        (x_5).value_write, value : (x_5).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_18).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (x_20).info_write, info : (x_20).info, value_write : (Bool)'(True),
        value : ((x_15).msg).value});
        let x_22 <- cache_00_writeRq(x_21);
        let x_23 <- releaseDL00((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_17)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_17)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_17)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h6),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        ((x_15).msg).value}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 = (wl00);
        when (! ((x_26).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_12;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((((x_10).dir_st) == ((Bit#(3))'(3'h1))) || ((((x_10).dir_st) ==
        ((Bit#(3))'(3'h2))) && (((x_10).dir_sharers) == (((Bit#(4))'(4'h1))
        << (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))), noAction);

        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_19 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_18)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_20 = (Struct3 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_19).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct3 x_21 = (Struct3 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_20).info).mesi_status, mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_00_writeRq(x_21);
        let x_23 <- releaseUL00((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_25 <- makeEnq_parentChildren00(x_24);
        let x_26 = (wl00);
        when (! ((x_26).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_13;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((Bool)'(True)) && ((!
        ((((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)})[1:0])))) ==
        ((Bit#(4))'(4'h0)))) && (((x_10).dir_st) == ((Bit#(3))'(3'h2)))))),
        noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = ((x_13).ul_msg);
        Bit#(4) x_17 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct3 x_18 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        let x_19 <- cache_00_writeRq(x_18);
        let x_20 <- transferUpDown00(Struct17 {r_dl_addr : (x_11).addr,
        r_dl_rss_from : ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) <<
        ((x_17)[1:0])))});
        let x_21 <- broadcast_parentChildren00(Struct13 {cs_inds :
        ((x_10).dir_sharers) & (~(((Bit#(4))'(4'h1)) << ((x_17)[1:0]))),
        cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ : (Bool)'(False), addr
        : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 = (wl00);
        when (! ((x_22).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_161;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'ha)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h4), dir_excl : (x_16)[1:0], dir_sharers :
        (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        let x_21 <- releaseDL00((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hb),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_170;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((x_10).dir_st) == ((Bit#(3))'(3'h1)), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct3 x_16 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_17 = (Struct3 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_171;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when ((! ((x_9) < ((Bit#(3))'(3'h3)))) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h1))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct3 x_16 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_17 = (Struct3 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_00_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren00(x_19);
        let x_21 = (wl00);
        when (! ((x_21).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_190;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_191;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && ((! (((x_10).dir_st) < ((Bit#(3))'(3'h3))))
        && (! (((Bit#(3))'(3'h4)) < ((x_10).dir_st)))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : ((Bit#(4))'(4'h0)) | (((Bit#(4))'(4'h1)) <<
        (({((Bit#(2))'(2'h1)),((x_10).dir_excl)})[1:0])), r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        Struct10 x_17 = (Struct10 {enq_type :
        ((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) :
        (((({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ({((Bit#(2))'(2'h2)),((x_10).dir_excl)})[1:0], enq_msg :
        Struct2 {id : (Bit#(6))'(6'he), type_ : (Bool)'(False), addr :
        (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 <- makeEnq_parentChildren00(x_17);
        let x_19 = (wl00);
        when (! ((x_19).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_192;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable00((x_11).addr);
        when (x_14, noAction);
        when (((Bool)'(True)) && (((Bool)'(True)) && (((x_10).dir_st) ==
        ((Bit#(3))'(3'h2)))), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- registerDL00(Struct12 {r_dl_rsb : (Bool)'(True), r_dl_msg
        : x_15, r_dl_rss_from : (x_10).dir_sharers, r_dl_rsbTo :
        (Bit#(4))'(4'h4)});
        let x_17 <- broadcast_parentChildren00(Struct13 {cs_inds :
        (x_10).dir_sharers, cs_msg : Struct2 {id : (Bit#(6))'(6'hc), type_ :
        (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_11010;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'hc)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        let x_21 <- releaseDL00((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hd),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_11011;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_3).rl_valid) && ((x_3).rl_line_valid), noAction);
        Struct3 x_4 = ((x_3).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_3).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        let x_13 <- downLockGet00((x_11).addr);
        when ((x_13).valid, noAction);
        Struct7 x_14 = ((x_13).data);
        when ((x_14).dl_valid, noAction);
        when ((x_14).dl_rsb, noAction);
        when ((((x_14).dl_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_14).dl_msg).id) == ((Bit#(6))'(6'he)), noAction);
        when (((x_14).dl_rss_recv) == ((x_14).dl_rss_from), noAction);
        when ((Bool)'(True), noAction);
        crsrl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = ((x_14).dl_msg);
        Bit#(4) x_16 = ((x_14).dl_rsbTo);
        Struct3 x_17 = (Struct3 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : ((x_5).info).mesi_status, mesi_dir_st : (Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_st, mesi_dir_sharers : (((Struct8 {dir_st :
        (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_st) == ((Bit#(3))'(3'h2)) ? ((Struct8 {dir_st
        : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers :
        (Bit#(4))'(4'h0)}).dir_sharers) : (((Bit#(4))'(4'h1)) << ((Struct8
        {dir_st : (Bit#(3))'(3'h1), dir_excl : (Bit#(2))'(2'h0), dir_sharers
        : (Bit#(4))'(4'h0)}).dir_excl)))}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct3 x_18 = (Struct3 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct3 x_19 = (Struct3 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_00_writeRq(x_19);
        let x_21 <- releaseDL00((x_11).addr);
        Struct10 x_22 = (Struct10 {enq_type : (((x_16)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_16)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_16)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'hf),
        type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_23 <- makeEnq_parentChildren00(x_22);
        let x_24 = (wl00);
        when (! ((x_24).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_00_20;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        let x_3 <- cache_00_getVictim();
        Struct3 x_4 = (Struct3 {addr : (x_3).addr, info_hit : (x_3).info_hit,
        info_way : (x_3).info_way, info_write : (x_3).info_write, info :
        Struct4 {mesi_owned : ((x_3).info).mesi_owned, mesi_status :
        ((((x_3).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable00((x_10).addr);
        when (x_13, noAction);
        when (((x_7) == ((Bool)'(False))) && (((((Bit#(3))'(3'h0)) < (x_8))
        && ((x_8) < ((Bit#(3))'(3'h4)))) && (((x_9).dir_st) ==
        ((Bit#(3))'(3'h1)))), noAction);
        let x_14 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_10).addr, value
        : (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_16 <- makeEnq_parentChildren00(x_15);
        let x_17 = (wl00);
        when (! ((x_17).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_21;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        let x_3 <- cache_00_getVictim();
        Struct3 x_4 = (Struct3 {addr : (x_3).addr, info_hit : (x_3).info_hit,
        info_way : (x_3).info_way, info_write : (x_3).info_write, info :
        Struct4 {mesi_owned : ((x_3).info).mesi_owned, mesi_status :
        ((((x_3).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable00((x_10).addr);
        when (x_13, noAction);
        when ((((x_9).dir_st) == ((Bit#(3))'(3'h1))) && ((((x_7) ==
        ((Bool)'(True))) && (((Bit#(3))'(3'h1)) < (x_8))) || (((x_7) ==
        ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) && ((x_8) <
        ((Bit#(3))'(3'h3)))))), noAction);
        let x_14 <- registerUL00(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_10).addr, value
        : x_5}});
        let x_16 <- makeEnq_parentChildren00(x_15);
        let x_17 = (wl00);
        when (! ((x_17).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_00_22;
        let x_0 = (rr00);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl00);
        let x_2 = (crqrl00);
        let x_3 = (crsrl00);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct3 x_4 = ((x_1).rl_line);
        Struct3 x_5 = (Struct3 {addr : (x_4).addr, info_hit : (x_4).info_hit,
        info_way : (x_4).info_way, info_write : (x_4).info_write, info :
        Struct4 {mesi_owned : ((x_4).info).mesi_owned, mesi_status :
        ((((x_4).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet00((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable00((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl00 <=
        (Struct1)'(Struct1 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL00((x_11).addr);
        let x_18 = (wl00);
        when (! ((x_18).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_00_removeVictim(x_19);
        let x_21 = (crqrl00);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl00 <= Struct1 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct3 {addr : x_19, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end
        let x_23 = (crsrl00);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl00 <= Struct1 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct3 {addr : x_19, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end

    endrule

    (* descending_urgency = "rule_00_23, rule_00_20, rule_00_21" *)
    rule rule_00_23;
        let x_0 = (prl00);
        let x_1 = (crqrl00);
        let x_2 = (crsrl00);
        let x_3 <- cache_00_getVictim();
        Struct3 x_4 = (Struct3 {addr : (x_3).addr, info_hit : (x_3).info_hit,
        info_way : (x_3).info_way, info_write : (x_3).info_write, info :
        Struct4 {mesi_owned : ((x_3).info).mesi_owned, mesi_status :
        ((((x_3).info).mesi_status) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        let x_13 <- upLockable00((x_10).addr);
        when (x_13, noAction);
        let x_14 <- downLockable00((x_10).addr);
        when (x_14, noAction);
        when ((((x_8) == ((Bit#(3))'(3'h1))) && (! (((x_9).dir_st) ==
        ((Bit#(3))'(3'h3))))) || (((x_8) == ((Bit#(3))'(3'h2))) && ((x_7) ==
        ((Bool)'(False)))), noAction);
        let x_15 = (wl00);
        when (! ((x_15).wl_valid), noAction);
        wl00 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_16 = ((x_10).addr);
        let x_17 <- cache_00_removeVictim(x_16);
        let x_18 = (crqrl00);
        if ((((x_18).rl_valid) && ((x_18).rl_line_valid)) &&
        ((((x_18).rl_msg).addr) == (x_16))) begin

            crqrl00 <= Struct1 {rl_valid : (x_18).rl_valid, rl_cmidx :
            (x_18).rl_cmidx, rl_msg : (x_18).rl_msg, rl_line_valid :
            (x_18).rl_line_valid, rl_line : Struct3 {addr : x_16, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end
        let x_20 = (crsrl00);
        if ((((x_20).rl_valid) && ((x_20).rl_line_valid)) &&
        ((((x_20).rl_msg).addr) == (x_16))) begin

            crsrl00 <= Struct1 {rl_valid : (x_20).rl_valid, rl_cmidx :
            (x_20).rl_cmidx, rl_msg : (x_20).rl_msg, rl_line_valid :
            (x_20).rl_line_valid, rl_line : Struct3 {addr : x_16, info_hit :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct3)'(Struct3 {addr: 64'h0, info_hit: False, info_way: 4'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end

    endrule

    rule rule_00_7890;
        let x_0 = (wl00);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl00 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_00_7891;
        let x_0 = (wl00);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_00_writeRs();
        let x_2 = (prl00);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl00);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl00);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl00 <= Struct1 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl00 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module74;
endinterface


module mkModule74#(function ActionValue#(Struct24) cache_000_writeRs(),
  function Action cache_000_removeVictim(Bit#(64) _),
  function ActionValue#(Struct24) cache_000_getVictim(),
  function Action releaseUL000(Bit#(64) _),
  function Action cache_000_writeRq(Struct24 _),
  function ActionValue#(Struct15) upLockGet000(Bit#(64) _),
  function Action registerUL000(Struct11 _),
  function ActionValue#(Bool) cache_000_hasVictimSlot(),
  function Action makeEnq_parentChildren000(Struct10 _),
  function ActionValue#(Bool) downLockable000(Bit#(64) _),
  function ActionValue#(Bool) upLockable000(Bit#(64) _),
  function ActionValue#(Struct24) cache_000_readRs(),
  function ActionValue#(Struct2) deq_fifo00000(),
  function ActionValue#(Struct6) downLockRssFull000(),
  function Action cache_000_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0002()) (Module74);
    Reg#(Bit#(1)) rr000 <- mkReg(unpack(0));
    Reg#(Struct23) prl000 <- mkReg(unpack(0));
    Reg#(Struct23) crqrl000 <- mkReg(unpack(0));
    Reg#(Struct23) crsrl000 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc000 <- mkReg(unpack(0));
    Reg#(Struct5) wl000 <- mkReg(unpack(0));

    rule rr_000;let x_0 = (rr000);
                rr000 <= (x_0) + ((Bit#(1))'(1'h1));

    endrule

    rule rule_000_1230;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo0002();
        prl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc000 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_000_readRq((x_3).addr);

    endrule

    rule rule_000_1232;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull000();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc000 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_000_readRq((x_4).addr);

    endrule

    rule rule_000_123100000;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00000();
        crqrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc000 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_000_readRq((x_3).addr);

    endrule

    rule rule_000_456;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        let x_3 <- cache_000_readRs();
        let x_4 = (rlc000);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl000 <= Struct23 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl000 <= Struct23 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl000 <= Struct23 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_000_00;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren000(x_17);
        let x_19 = (wl000);
        when (! ((x_19).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_01;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_020;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_000_writeRq(x_20);
        let x_22 <- releaseUL000((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren000(x_23);
        let x_25 = (wl000);
        when (! ((x_25).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_021;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_000_writeRq(x_20);
        let x_22 <- releaseUL000((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren000(x_23);
        let x_25 = (wl000);
        when (! ((x_25).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_03;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_100;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_000_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren000(x_21);
        let x_23 = (wl000);
        when (! ((x_23).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_101;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_11;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable000((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_000_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren000(x_18);
        let x_20 = (wl000);
        when (! ((x_20).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_12;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_000_writeRq(x_21);
        let x_23 <- releaseUL000((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_25 <- makeEnq_parentChildren000(x_24);
        let x_26 = (wl000);
        when (! ((x_26).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_130;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_131;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable000((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_000_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h4))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h4))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h4))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren000(x_19);
        let x_21 = (wl000);
        when (! ((x_21).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_000_20;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        let x_3 <- cache_000_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable000((x_10).addr);
        when (x_13, noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        let x_14 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_10).addr, value
        : (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_16 <- makeEnq_parentChildren000(x_15);
        let x_17 = (wl000);
        when (! ((x_17).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_000_20, rule_000_21" *)
    rule rule_000_21;
        let x_0 = (prl000);
        let x_1 = (crqrl000);
        let x_2 = (crsrl000);
        let x_3 <- cache_000_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable000((x_10).addr);
        when (x_13, noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        let x_14 <- registerUL000(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h0))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h0))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h0))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_10).addr, value
        : x_5}});
        let x_16 <- makeEnq_parentChildren000(x_15);
        let x_17 = (wl000);
        when (! ((x_17).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_000_22;
        let x_0 = (rr000);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl000);
        let x_2 = (crqrl000);
        let x_3 = (crsrl000);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet000((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable000((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl000 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL000((x_11).addr);
        let x_18 = (wl000);
        when (! ((x_18).wl_valid), noAction);
        wl000 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_000_removeVictim(x_19);
        let x_21 = (crqrl000);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl000 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end
        let x_23 = (crsrl000);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl000 <= Struct23 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end

    endrule

    rule rule_000_7890;
        let x_0 = (wl000);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl000 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_000_7891;
        let x_0 = (wl000);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_000_writeRs();
        let x_2 = (prl000);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl000);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl000);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl000 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl000 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module75;
endinterface


module mkModule75#(function ActionValue#(Struct24) cache_001_writeRs(),
  function Action cache_001_removeVictim(Bit#(64) _),
  function ActionValue#(Struct24) cache_001_getVictim(),
  function Action releaseUL001(Bit#(64) _),
  function Action cache_001_writeRq(Struct24 _),
  function ActionValue#(Struct15) upLockGet001(Bit#(64) _),
  function Action registerUL001(Struct11 _),
  function ActionValue#(Bool) cache_001_hasVictimSlot(),
  function Action makeEnq_parentChildren001(Struct10 _),
  function ActionValue#(Bool) downLockable001(Bit#(64) _),
  function ActionValue#(Bool) upLockable001(Bit#(64) _),
  function ActionValue#(Struct24) cache_001_readRs(),
  function ActionValue#(Struct2) deq_fifo00100(),
  function ActionValue#(Struct6) downLockRssFull001(),
  function Action cache_001_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0012()) (Module75);
    Reg#(Bit#(1)) rr001 <- mkReg(unpack(0));
    Reg#(Struct23) prl001 <- mkReg(unpack(0));
    Reg#(Struct23) crqrl001 <- mkReg(unpack(0));
    Reg#(Struct23) crsrl001 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc001 <- mkReg(unpack(0));
    Reg#(Struct5) wl001 <- mkReg(unpack(0));

    rule rr_001;let x_0 = (rr001);
                rr001 <= (x_0) + ((Bit#(1))'(1'h1));

    endrule

    rule rule_001_1230;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo0012();
        prl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc001 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_001_readRq((x_3).addr);

    endrule

    rule rule_001_1232;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull001();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc001 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_001_readRq((x_4).addr);

    endrule

    rule rule_001_123100100;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00100();
        crqrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc001 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_001_readRq((x_3).addr);

    endrule

    rule rule_001_456;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        let x_3 <- cache_001_readRs();
        let x_4 = (rlc001);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl001 <= Struct23 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl001 <= Struct23 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl001 <= Struct23 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_001_00;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren001(x_17);
        let x_19 = (wl001);
        when (! ((x_19).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_01;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_020;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_001_writeRq(x_20);
        let x_22 <- releaseUL001((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren001(x_23);
        let x_25 = (wl001);
        when (! ((x_25).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_021;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_001_writeRq(x_20);
        let x_22 <- releaseUL001((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren001(x_23);
        let x_25 = (wl001);
        when (! ((x_25).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_03;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_100;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_001_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren001(x_21);
        let x_23 = (wl001);
        when (! ((x_23).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_101;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_11;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable001((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_001_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren001(x_18);
        let x_20 = (wl001);
        when (! ((x_20).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_12;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_001_writeRq(x_21);
        let x_23 <- releaseUL001((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_25 <- makeEnq_parentChildren001(x_24);
        let x_26 = (wl001);
        when (! ((x_26).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_130;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_131;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable001((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_001_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h5))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h5))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h5))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren001(x_19);
        let x_21 = (wl001);
        when (! ((x_21).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_001_20;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        let x_3 <- cache_001_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable001((x_10).addr);
        when (x_13, noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        let x_14 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_10).addr, value
        : (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_16 <- makeEnq_parentChildren001(x_15);
        let x_17 = (wl001);
        when (! ((x_17).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_001_20, rule_001_21" *)
    rule rule_001_21;
        let x_0 = (prl001);
        let x_1 = (crqrl001);
        let x_2 = (crsrl001);
        let x_3 <- cache_001_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable001((x_10).addr);
        when (x_13, noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        let x_14 <- registerUL001(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h1))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h1))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h1))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_10).addr, value
        : x_5}});
        let x_16 <- makeEnq_parentChildren001(x_15);
        let x_17 = (wl001);
        when (! ((x_17).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_001_22;
        let x_0 = (rr001);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl001);
        let x_2 = (crqrl001);
        let x_3 = (crsrl001);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet001((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable001((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl001 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL001((x_11).addr);
        let x_18 = (wl001);
        when (! ((x_18).wl_valid), noAction);
        wl001 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_001_removeVictim(x_19);
        let x_21 = (crqrl001);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl001 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end
        let x_23 = (crsrl001);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl001 <= Struct23 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end

    endrule

    rule rule_001_7890;
        let x_0 = (wl001);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl001 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_001_7891;
        let x_0 = (wl001);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_001_writeRs();
        let x_2 = (prl001);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl001);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl001);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl001 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl001 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module76;
endinterface


module mkModule76#(function ActionValue#(Struct24) cache_002_writeRs(),
  function Action cache_002_removeVictim(Bit#(64) _),
  function ActionValue#(Struct24) cache_002_getVictim(),
  function Action releaseUL002(Bit#(64) _),
  function Action cache_002_writeRq(Struct24 _),
  function ActionValue#(Struct15) upLockGet002(Bit#(64) _),
  function Action registerUL002(Struct11 _),
  function ActionValue#(Bool) cache_002_hasVictimSlot(),
  function Action makeEnq_parentChildren002(Struct10 _),
  function ActionValue#(Bool) downLockable002(Bit#(64) _),
  function ActionValue#(Bool) upLockable002(Bit#(64) _),
  function ActionValue#(Struct24) cache_002_readRs(),
  function ActionValue#(Struct2) deq_fifo00200(),
  function ActionValue#(Struct6) downLockRssFull002(),
  function Action cache_002_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0022()) (Module76);
    Reg#(Bit#(1)) rr002 <- mkReg(unpack(0));
    Reg#(Struct23) prl002 <- mkReg(unpack(0));
    Reg#(Struct23) crqrl002 <- mkReg(unpack(0));
    Reg#(Struct23) crsrl002 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc002 <- mkReg(unpack(0));
    Reg#(Struct5) wl002 <- mkReg(unpack(0));

    rule rr_002;let x_0 = (rr002);
                rr002 <= (x_0) + ((Bit#(1))'(1'h1));

    endrule

    rule rule_002_1230;
        let x_0 = (prl002);
        let x_1 = (crqrl002);
        let x_2 = (crsrl002);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo0022();
        prl002 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc002 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_002_readRq((x_3).addr);

    endrule

    rule rule_002_1232;
        let x_0 = (prl002);
        let x_1 = (crqrl002);
        let x_2 = (crsrl002);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull002();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl002 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc002 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_002_readRq((x_4).addr);

    endrule

    rule rule_002_123100200;
        let x_0 = (prl002);
        let x_1 = (crqrl002);
        let x_2 = (crsrl002);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00200();
        crqrl002 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc002 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_002_readRq((x_3).addr);

    endrule

    rule rule_002_456;
        let x_0 = (prl002);
        let x_1 = (crqrl002);
        let x_2 = (crsrl002);
        let x_3 <- cache_002_readRs();
        let x_4 = (rlc002);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl002 <= Struct23 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl002 <= Struct23 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl002 <= Struct23 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_002_00;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable002((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable002((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren002(x_17);
        let x_19 = (wl002);
        when (! ((x_19).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_002_01;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable002((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_002_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL002(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren002(x_18);
        let x_20 = (wl002);
        when (! ((x_20).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_002_020;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_002_writeRq(x_20);
        let x_22 <- releaseUL002((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren002(x_23);
        let x_25 = (wl002);
        when (! ((x_25).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_021;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_002_writeRq(x_20);
        let x_22 <- releaseUL002((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren002(x_23);
        let x_25 = (wl002);
        when (! ((x_25).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_03;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable002((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren002(x_19);
        let x_21 = (wl002);
        when (! ((x_21).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_100;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable002((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable002((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_002_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren002(x_21);
        let x_23 = (wl002);
        when (! ((x_23).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_101;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable002((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable002((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren002(x_19);
        let x_21 = (wl002);
        when (! ((x_21).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_11;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable002((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_002_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL002(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren002(x_18);
        let x_20 = (wl002);
        when (! ((x_20).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_002_12;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_002_writeRq(x_21);
        let x_23 <- releaseUL002((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_25 <- makeEnq_parentChildren002(x_24);
        let x_26 = (wl002);
        when (! ((x_26).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_130;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable002((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren002(x_19);
        let x_21 = (wl002);
        when (! ((x_21).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_131;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable002((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_002_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h6))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h6))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h6))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren002(x_19);
        let x_21 = (wl002);
        when (! ((x_21).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_002_20;
        let x_0 = (prl002);
        let x_1 = (crqrl002);
        let x_2 = (crsrl002);
        let x_3 <- cache_002_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable002((x_10).addr);
        when (x_13, noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        let x_14 <- registerUL002(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_10).addr, value
        : (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_16 <- makeEnq_parentChildren002(x_15);
        let x_17 = (wl002);
        when (! ((x_17).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_002_20, rule_002_21" *)
    rule rule_002_21;
        let x_0 = (prl002);
        let x_1 = (crqrl002);
        let x_2 = (crsrl002);
        let x_3 <- cache_002_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable002((x_10).addr);
        when (x_13, noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        let x_14 <- registerUL002(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h2))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h2))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h2))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_10).addr, value
        : x_5}});
        let x_16 <- makeEnq_parentChildren002(x_15);
        let x_17 = (wl002);
        when (! ((x_17).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_002_22;
        let x_0 = (rr002);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl002);
        let x_2 = (crqrl002);
        let x_3 = (crsrl002);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet002((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable002((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl002 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL002((x_11).addr);
        let x_18 = (wl002);
        when (! ((x_18).wl_valid), noAction);
        wl002 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_002_removeVictim(x_19);
        let x_21 = (crqrl002);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl002 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end
        let x_23 = (crsrl002);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl002 <= Struct23 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end

    endrule

    rule rule_002_7890;
        let x_0 = (wl002);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl002 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_002_7891;
        let x_0 = (wl002);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_002_writeRs();
        let x_2 = (prl002);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl002 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl002);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl002 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl002);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl002 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl002 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule

interface Module77;
endinterface


module mkModule77#(function ActionValue#(Struct24) cache_003_writeRs(),
  function Action cache_003_removeVictim(Bit#(64) _),
  function ActionValue#(Struct24) cache_003_getVictim(),
  function Action releaseUL003(Bit#(64) _),
  function Action cache_003_writeRq(Struct24 _),
  function ActionValue#(Struct15) upLockGet003(Bit#(64) _),
  function Action registerUL003(Struct11 _),
  function ActionValue#(Bool) cache_003_hasVictimSlot(),
  function Action makeEnq_parentChildren003(Struct10 _),
  function ActionValue#(Bool) downLockable003(Bit#(64) _),
  function ActionValue#(Bool) upLockable003(Bit#(64) _),
  function ActionValue#(Struct24) cache_003_readRs(),
  function ActionValue#(Struct2) deq_fifo00300(),
  function ActionValue#(Struct6) downLockRssFull003(),
  function Action cache_003_readRq(Bit#(64) _),
  function ActionValue#(Struct2) deq_fifo0032()) (Module77);
    Reg#(Bit#(1)) rr003 <- mkReg(unpack(0));
    Reg#(Struct23) prl003 <- mkReg(unpack(0));
    Reg#(Struct23) crqrl003 <- mkReg(unpack(0));
    Reg#(Struct23) crsrl003 <- mkReg(unpack(0));
    Reg#(Bit#(2)) rlc003 <- mkReg(unpack(0));
    Reg#(Struct5) wl003 <- mkReg(unpack(0));

    rule rr_003;let x_0 = (rr003);
                rr003 <= (x_0) + ((Bit#(1))'(1'h1));

    endrule

    rule rule_003_1230;
        let x_0 = (prl003);
        let x_1 = (crqrl003);
        let x_2 = (crsrl003);
        when (! ((x_0).rl_valid), noAction);
        let x_3 <- deq_fifo0032();
        prl003 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc003 <= (Bit#(2))'(2'h2);
        let x_4 <- cache_003_readRq((x_3).addr);

    endrule

    rule rule_003_1232;
        let x_0 = (prl003);
        let x_1 = (crqrl003);
        let x_2 = (crsrl003);
        when (! ((x_2).rl_valid), noAction);
        let x_3 <- downLockRssFull003();
        when ((x_3).valid, noAction);
        Struct2 x_4 = (((x_3).data).dl_msg);
        crsrl003 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_4, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc003 <= (Bit#(2))'(2'h1);
        let x_5 <- cache_003_readRq((x_4).addr);

    endrule

    rule rule_003_123100300;
        let x_0 = (prl003);
        let x_1 = (crqrl003);
        let x_2 = (crsrl003);
        when (! ((x_1).rl_valid), noAction);
        let x_3 <- deq_fifo00300();
        crqrl003 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
        (Bit#(2))'(2'h0), rl_msg : x_3, rl_line_valid : (Bool)'(False),
        rl_line :
        (Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})};

        rlc003 <= (Bit#(2))'(2'h0);
        let x_4 <- cache_003_readRq((x_3).addr);

    endrule

    rule rule_003_456;
        let x_0 = (prl003);
        let x_1 = (crqrl003);
        let x_2 = (crsrl003);
        let x_3 <- cache_003_readRs();
        let x_4 = (rlc003);
        if ((x_4) == ((Bit#(2))'(2'h0))) begin

            crqrl003 <= Struct23 {rl_valid : (x_1).rl_valid, rl_cmidx :
            (x_1).rl_cmidx, rl_msg : (x_1).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_3};

        end else begin

            if ((x_4) == ((Bit#(2))'(2'h1))) begin

                crsrl003 <= Struct23 {rl_valid : (x_2).rl_valid, rl_cmidx :
                (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end else begin

                prl003 <= Struct23 {rl_valid : (x_0).rl_valid, rl_cmidx :
                (x_0).rl_cmidx, rl_msg : (x_0).rl_msg, rl_line_valid :
                (Bool)'(True), rl_line : x_3};

            end

        end

    endrule

    rule rule_003_00;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable003((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable003((x_11).addr);
        when (x_15, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        crqrl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct10 x_17 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h1), type_ : (Bool)'(True), addr : (x_16).addr, value :
        x_6}});
        let x_18 <- makeEnq_parentChildren003(x_17);
        let x_19 = (wl003);
        when (! ((x_19).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_003_01;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h0)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable003((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h1)) < (x_9)), noAction);
        crqrl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_003_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL003(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h2), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren003(x_18);
        let x_20 = (wl003);
        when (! ((x_20).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_003_020;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h3)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_003_writeRq(x_20);
        let x_22 <- releaseUL003((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren003(x_23);
        let x_25 = (wl003);
        when (! ((x_25).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_021;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h4)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h0)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h3), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (x_19).info_write, info : (x_19).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_21 <- cache_003_writeRq(x_20);
        let x_22 <- releaseUL003((x_11).addr);
        Struct10 x_23 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h1),
        type_ : (Bool)'(True), addr : (x_16).addr, value : (x_16).value}});

        let x_24 <- makeEnq_parentChildren003(x_23);
        let x_25 = (wl003);
        when (! ((x_25).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_03;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h5)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable003((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h2))), noAction);
        prl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h2), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h6), type_ : (Bool)'(True), addr : (x_15).addr, value :
        x_6}});
        let x_20 <- makeEnq_parentChildren003(x_19);
        let x_21 = (wl003);
        when (! ((x_21).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_100;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable003((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable003((x_11).addr);
        when (x_15, noAction);
        when ((x_9) == ((Bit#(3))'(3'h3)), noAction);
        crqrl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        Struct24 x_18 = (Struct24 {addr : (x_17).addr, info_hit :
        (x_17).info_hit, info_way : (x_17).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_17).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_17).info).mesi_dir_st, mesi_dir_sharers :
        ((x_17).info).mesi_dir_sharers}, value_write : (x_17).value_write,
        value : (x_17).value});
        Struct24 x_19 = (Struct24 {addr : (x_18).addr, info_hit :
        (x_18).info_hit, info_way : (x_18).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_18).info).mesi_status, mesi_dir_st :
        ((x_18).info).mesi_dir_st, mesi_dir_sharers :
        ((x_18).info).mesi_dir_sharers}, value_write : (x_18).value_write,
        value : (x_18).value});
        let x_20 <- cache_003_writeRq(x_19);
        Struct10 x_21 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_22 <- makeEnq_parentChildren003(x_21);
        let x_23 = (wl003);
        when (! ((x_23).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_101;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable003((x_11).addr);
        when (x_14, noAction);
        let x_15 <- downLockable003((x_11).addr);
        when (x_15, noAction);
        when (((x_8) == ((Bool)'(True))) && ((x_9) == ((Bit#(3))'(3'h4))),
        noAction);
        crqrl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct24 x_17 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_16).value});
        let x_18 <- cache_003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h8))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h8))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h8))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h9), type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren003(x_19);
        let x_21 = (wl003);
        when (! ((x_21).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_11;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h1)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_2).rl_valid) && ((x_2).rl_line_valid), noAction);
        when (((x_2).rl_cmidx) == ((Bit#(2))'(2'h0)), noAction);
        Struct24 x_4 = ((x_2).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_2).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h8)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- upLockable003((x_11).addr);
        when (x_14, noAction);
        when (! (((Bit#(3))'(3'h2)) < (x_9)), noAction);
        crqrl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        let x_16 <- cache_003_hasVictimSlot();
        when (! (x_16), noAction);
        let x_17 <- registerUL003(Struct11 {r_ul_rsb : (Bool)'(True),
        r_ul_msg : x_15, r_ul_rsbTo : ((Bit#(4))'(4'h8))[1:0]});
        Struct10 x_18 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'ha), type_ : (Bool)'(False), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_19 <- makeEnq_parentChildren003(x_18);
        let x_20 = (wl003);
        when (! ((x_20).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_003_12;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hb)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((((x_13).ul_msg).type_) == ((Bool)'(False)), noAction);
        when ((((x_13).ul_msg).id) == ((Bit#(6))'(6'h8)), noAction);
        when ((x_13).ul_valid, noAction);
        when ((x_13).ul_rsb, noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        Struct2 x_17 = ((x_13).ul_msg);
        Bit#(4) x_18 = ({((Bit#(2))'(2'h2)),((x_13).ul_rsbTo)});
        Struct24 x_19 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (x_5).info_write, info : (x_5).info, value_write : (Bool)'(True),
        value : (x_17).value});
        Struct24 x_20 = (Struct24 {addr : (x_19).addr, info_hit :
        (x_19).info_hit, info_way : (x_19).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(True),
        mesi_status : ((x_19).info).mesi_status, mesi_dir_st :
        ((x_19).info).mesi_dir_st, mesi_dir_sharers :
        ((x_19).info).mesi_dir_sharers}, value_write : (x_19).value_write,
        value : (x_19).value});
        Struct24 x_21 = (Struct24 {addr : (x_20).addr, info_hit :
        (x_20).info_hit, info_way : (x_20).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_20).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h4), mesi_dir_st :
        ((x_20).info).mesi_dir_st, mesi_dir_sharers :
        ((x_20).info).mesi_dir_sharers}, value_write : (x_20).value_write,
        value : (x_20).value});
        let x_22 <- cache_003_writeRq(x_21);
        let x_23 <- releaseUL003((x_11).addr);
        Struct10 x_24 = (Struct10 {enq_type : (((x_18)[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : ((((x_18)[3:2]) ==
        ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : (x_18)[1:0], enq_msg : Struct2 {id : (Bit#(6))'(6'h9),
        type_ : (Bool)'(True), addr : (x_16).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_25 <- makeEnq_parentChildren003(x_24);
        let x_26 = (wl003);
        when (! ((x_26).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_130;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'hc)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable003((x_11).addr);
        when (x_14, noAction);
        when ((Bool)'(True), noAction);
        prl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hd), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren003(x_19);
        let x_21 = (wl003);
        when (! ((x_21).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_131;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        Struct9 x_12 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_13 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'he)), noAction);
        when (! ((x_11).type_), noAction);
        let x_14 <- downLockable003((x_11).addr);
        when (x_14, noAction);
        when (! ((x_9) < ((Bit#(3))'(3'h3))), noAction);
        prl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_15 = (x_11);
        Struct24 x_16 = (Struct24 {addr : (x_5).addr, info_hit :
        (x_5).info_hit, info_way : (x_5).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : ((x_5).info).mesi_owned,
        mesi_status : (Bit#(3))'(3'h1), mesi_dir_st :
        ((x_5).info).mesi_dir_st, mesi_dir_sharers :
        ((x_5).info).mesi_dir_sharers}, value_write : (x_5).value_write,
        value : (x_5).value});
        Struct24 x_17 = (Struct24 {addr : (x_16).addr, info_hit :
        (x_16).info_hit, info_way : (x_16).info_way, info_write :
        (Bool)'(True), info : Struct4 {mesi_owned : (Bool)'(False),
        mesi_status : ((x_16).info).mesi_status, mesi_dir_st :
        ((x_16).info).mesi_dir_st, mesi_dir_sharers :
        ((x_16).info).mesi_dir_sharers}, value_write : (x_16).value_write,
        value : (x_16).value});
        let x_18 <- cache_003_writeRq(x_17);
        Struct10 x_19 = (Struct10 {enq_type : ((((Bit#(4))'(4'h7))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h7))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h7))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'hf), type_ : (Bool)'(True), addr : (x_15).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_20 <- makeEnq_parentChildren003(x_19);
        let x_21 = (wl003);
        when (! ((x_21).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(True)};

    endrule

    rule rule_003_20;
        let x_0 = (prl003);
        let x_1 = (crqrl003);
        let x_2 = (crsrl003);
        let x_3 <- cache_003_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable003((x_10).addr);
        when (x_13, noAction);
        when (((x_7) == ((Bool)'(False))) && ((((Bit#(3))'(3'h0)) < (x_8)) &&
        ((x_8) < ((Bit#(3))'(3'h4)))), noAction);
        let x_14 <- registerUL003(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h14), type_ : (Bool)'(False), addr : (x_10).addr, value
        : (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))}});
        let x_16 <- makeEnq_parentChildren003(x_15);
        let x_17 = (wl003);
        when (! ((x_17).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    (* descending_urgency = "rule_003_20, rule_003_21" *)
    rule rule_003_21;
        let x_0 = (prl003);
        let x_1 = (crqrl003);
        let x_2 = (crsrl003);
        let x_3 <- cache_003_getVictim();
        Struct24 x_4 = (Struct24 {addr : (x_3).addr, info_hit :
        (x_3).info_hit, info_way : (x_3).info_way, info_write :
        (x_3).info_write, info : Struct4 {mesi_owned :
        ((x_3).info).mesi_owned, mesi_status : ((((x_3).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_3).info).mesi_status)), mesi_dir_st :
        ((((x_3).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_3).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_3).info).mesi_dir_sharers}, value_write : (x_3).value_write,
        value : (x_3).value});
        Vector#(4, Bit#(64)) x_5 = ((x_4).value);
        Struct4 x_6 = ((x_4).info);
        Bool x_7 = ((x_6).mesi_owned);
        Bit#(3) x_8 = ((x_6).mesi_status);
        Struct8 x_9 = (Struct8 {dir_st : (x_6).mesi_dir_st, dir_excl :
        ((((x_6).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_6).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_6).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_6).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_6).mesi_dir_sharers});
        Struct2 x_10 = (Struct2 {id : (Bit#(6))'(6'h0), type_ :
        (Bool)'(False), addr : (x_4).addr, value :
        (Vector#(4, Bit#(64)))'(vec(64'h0, 64'h0, 64'h0, 64'h0))});
        Struct9 x_11 =
        ((Struct9)'(Struct9 {ul_valid: False, ul_rsb: False, ul_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, ul_rsbTo: 2'h0}));

        Struct7 x_12 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (! ((x_10).type_), noAction);
        let x_13 <- upLockable003((x_10).addr);
        when (x_13, noAction);
        when (((Bit#(3))'(3'h0)) < (x_8), noAction);
        let x_14 <- registerUL003(Struct11 {r_ul_rsb : (Bool)'(False),
        r_ul_msg : x_10, r_ul_rsbTo : (Bit#(2))'(2'h0)});
        Struct10 x_15 = (Struct10 {enq_type : ((((Bit#(4))'(4'h3))[3:2]) ==
        ((Bit#(2))'(2'h2)) ? ((Bit#(2))'(2'h2)) : (((((Bit#(4))'(4'h3))[3:2])
        == ((Bit#(2))'(2'h0)) ? ((Bit#(2))'(2'h0)) : ((Bit#(2))'(2'h1))))),
        enq_ch_idx : ((Bit#(4))'(4'h3))[1:0], enq_msg : Struct2 {id :
        (Bit#(6))'(6'h15), type_ : (Bool)'(False), addr : (x_10).addr, value
        : x_5}});
        let x_16 <- makeEnq_parentChildren003(x_15);
        let x_17 = (wl003);
        when (! ((x_17).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};

    endrule

    rule rule_003_22;
        let x_0 = (rr003);
        when ((x_0) == ((Bit#(1))'(1'h0)), noAction);
        let x_1 = (prl003);
        let x_2 = (crqrl003);
        let x_3 = (crsrl003);
        when (((x_1).rl_valid) && ((x_1).rl_line_valid), noAction);
        Struct24 x_4 = ((x_1).rl_line);
        Struct24 x_5 = (Struct24 {addr : (x_4).addr, info_hit :
        (x_4).info_hit, info_way : (x_4).info_way, info_write :
        (x_4).info_write, info : Struct4 {mesi_owned :
        ((x_4).info).mesi_owned, mesi_status : ((((x_4).info).mesi_status) ==
        ((Bit#(3))'(3'h0)) ? ((Bit#(3))'(3'h1)) :
        (((x_4).info).mesi_status)), mesi_dir_st :
        ((((x_4).info).mesi_dir_st) == ((Bit#(3))'(3'h0)) ?
        ((Bit#(3))'(3'h1)) : (((x_4).info).mesi_dir_st)), mesi_dir_sharers :
        ((x_4).info).mesi_dir_sharers}, value_write : (x_4).value_write,
        value : (x_4).value});
        Vector#(4, Bit#(64)) x_6 = ((x_5).value);
        Struct4 x_7 = ((x_5).info);
        Bool x_8 = ((x_7).mesi_owned);
        Bit#(3) x_9 = ((x_7).mesi_status);
        Struct8 x_10 = (Struct8 {dir_st : (x_7).mesi_dir_st, dir_excl :
        ((((x_7).mesi_dir_sharers)[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((x_7).mesi_dir_sharers)[3:1])[0:0]) == ((Bit#(1))'(1'h1)) ?
        ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        (((((((x_7).mesi_dir_sharers)[3:1])[2:1])[0:0]) == ((Bit#(1))'(1'h1))
        ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((((((((x_7).mesi_dir_sharers)[3:1])[2:1])[1:1])[0:0]) ==
        ((Bit#(1))'(1'h1)) ? ((Bit#(2))'(2'h0)) : (((Bit#(2))'(2'h1)) +
        ((Bit#(2))'(2'h0))))))))))))), dir_sharers :
        (x_7).mesi_dir_sharers});
        Struct2 x_11 = ((x_1).rl_msg);
        let x_12 <- upLockGet003((x_11).addr);
        when ((x_12).valid, noAction);
        Struct9 x_13 = ((x_12).data);
        Struct7 x_14 =
        ((Struct7)'(Struct7 {dl_valid: False, dl_rsb: False, dl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, dl_rss_from: 4'h0, dl_rss_recv: 4'h0, dl_rss: vec(Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}), dl_rsbTo: 4'h0}));

        when (((x_11).id) == ((Bit#(6))'(6'h16)), noAction);
        when ((x_13).ul_valid, noAction);
        when (! ((x_13).ul_rsb), noAction);
        when ((x_11).type_, noAction);
        let x_15 <- downLockable003((x_11).addr);
        when (x_15, noAction);
        when ((Bool)'(True), noAction);
        prl003 <=
        (Struct23)'(Struct23 {rl_valid: False, rl_cmidx: 2'h0, rl_msg: Struct2 {id: 6'h0, type_: False, addr: 64'h0, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}, rl_line_valid: False, rl_line: Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)}});

        Struct2 x_16 = (x_11);
        let x_17 <- releaseUL003((x_11).addr);
        let x_18 = (wl003);
        when (! ((x_18).wl_valid), noAction);
        wl003 <= Struct5 {wl_valid : (Bool)'(True), wl_write_rq :
        (Bool)'(False)};
        Bit#(64) x_19 = ((x_11).addr);
        let x_20 <- cache_003_removeVictim(x_19);
        let x_21 = (crqrl003);
        if ((((x_21).rl_valid) && ((x_21).rl_line_valid)) &&
        ((((x_21).rl_msg).addr) == (x_19))) begin

            crqrl003 <= Struct23 {rl_valid : (x_21).rl_valid, rl_cmidx :
            (x_21).rl_cmidx, rl_msg : (x_21).rl_msg, rl_line_valid :
            (x_21).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end
        let x_23 = (crsrl003);
        if ((((x_23).rl_valid) && ((x_23).rl_line_valid)) &&
        ((((x_23).rl_msg).addr) == (x_19))) begin

            crsrl003 <= Struct23 {rl_valid : (x_23).rl_valid, rl_cmidx :
            (x_23).rl_cmidx, rl_msg : (x_23).rl_msg, rl_line_valid :
            (x_23).rl_line_valid, rl_line : Struct24 {addr : x_19, info_hit :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_hit,
            info_way :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_way,
            info_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info_write,
            info :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).info,
            value_write :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value_write,
            value :
            ((Struct24)'(Struct24 {addr: 64'h0, info_hit: False, info_way: 2'h0, info_write: False, info: Struct4 {mesi_owned: False, mesi_status: 3'h0, mesi_dir_st: 3'h0, mesi_dir_sharers: 4'h0}, value_write: False, value: vec(64'h0, 64'h0, 64'h0, 64'h0)})).value}};


        end else begin

        end

    endrule

    rule rule_003_7890;
        let x_0 = (wl003);
        when (((x_0).wl_valid) && (! ((x_0).wl_write_rq)), noAction);
        wl003 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    rule rule_003_7891;
        let x_0 = (wl003);
        when (((x_0).wl_valid) && ((x_0).wl_write_rq), noAction);
        let x_1 <- cache_003_writeRs();
        let x_2 = (prl003);
        if ((((x_2).rl_valid) && ((x_2).rl_line_valid)) &&
        ((((x_2).rl_msg).addr) == ((x_1).addr))) begin

            prl003 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_2).rl_cmidx, rl_msg : (x_2).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_4 = (crqrl003);
        if ((((x_4).rl_valid) && ((x_4).rl_line_valid)) &&
        ((((x_4).rl_msg).addr) == ((x_1).addr))) begin

            crqrl003 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_4).rl_cmidx, rl_msg : (x_4).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        let x_6 = (crsrl003);
        if ((((x_6).rl_valid) && ((x_6).rl_line_valid)) &&
        ((((x_6).rl_msg).addr) == ((x_1).addr))) begin

            crsrl003 <= Struct23 {rl_valid : (Bool)'(True), rl_cmidx :
            (x_6).rl_cmidx, rl_msg : (x_6).rl_msg, rl_line_valid :
            (Bool)'(True), rl_line : x_1};

        end else begin

        end
        wl003 <= (Struct5)'(Struct5 {wl_valid: False, wl_write_rq: False});

    endrule

    // No methods in this module
endmodule


// The CC interface is defined in the header part (thus in Header.bsv)

module mkCC#(function ActionValue#(Struct2) deq_fifo002(),
  function Action enq_fifo001(Struct2 _),
  function Action enq_fifo000(Struct2 _)) (CC);
    Module1 m1 <- mkModule1 ();
    Module2 m2 <- mkModule2 ();
    Module3 m3 <- mkModule3 ();
    Module4 m4 <- mkModule4 ();
    Module5 m5 <- mkModule5 ();
    Module6 m6 <- mkModule6 ();
    Module7 m7 <- mkModule7 ();
    Module8 m8 <- mkModule8 ();
    Module9 m9 <- mkModule9 ();
    Module10 m10 <- mkModule10 ();
    Module11 m11 <- mkModule11 ();
    Module12 m12 <- mkModule12 ();
    Module13 m13 <- mkModule13 ();
    Module14 m14 <- mkModule14 ();
    Module15 m15 <- mkModule15 ();
    Module16 m16 <- mkModule16 ();
    Module17 m17 <- mkModule17 ();
    Module18 m18 <- mkModule18 ();
    Module19 m19 <- mkModule19 ();
    Module20 m20 <- mkModule20 ();
    Module21 m21 <- mkModule21 ();
    Module22 m22 <- mkModule22 ();
    Module23 m23 <- mkModule23 ();
    Module24 m24 <- mkModule24 ();
    Module25 m25 <- mkModule25 ();
    Module26 m26 <- mkModule26 ();
    Module27 m27 <- mkModule27 ();
    Module28 m28 <- mkModule28 ();
    Module29 m29 <- mkModule29 ();
    Module30 m30 <- mkModule30 ();
    Module31 m31 <- mkModule31 ();
    Module32 m32 <- mkModule32 ();
    Module33 m33 <- mkModule33 ();
    Module34 m34 <- mkModule34 ();
    Module35 m35 <- mkModule35 ();
    Module36 m36 <- mkModule36 ();
    Module37 m37 <- mkModule37 ();
    Module38 m38 <- mkModule38 ();
    Module39 m39 <- mkModule39 ();
    Module40 m40 <- mkModule40 ();
    Module41 m41 <- mkModule41 ();
    Module42 m42 <- mkModule42 ();
    Module43 m43 <- mkModule43 ();
    Module44 m44 <- mkModule44 ();
    Module45 m45 <- mkModule45 ();
    Module46 m46 <- mkModule46 ();
    Module47 m47 <- mkModule47 ();
    Module48 m48 <- mkModule48 ();
    Module49 m49 <- mkModule49 ();
    Module50 m50 <- mkModule50 ();
    Module51 m51 <- mkModule51 ();
    Module52 m52 <- mkModule52 ();
    Module53 m53 <- mkModule53 ();
    Module54 m54 <- mkModule54 ();
    Module55 m55 <- mkModule55 ();
    Module56 m56 <- mkModule56 ();
    Module57 m57 <- mkModule57 ();
    Module58 m58 <- mkModule58 ();
    Module59 m59 <- mkModule59 ();
    Module60 m60 <- mkModule60 ();
    Module61 m61 <- mkModule61 ();
    Module62 m62 <- mkModule62 ();
    Module63 m63 <- mkModule63 (m1.putRq_infoRam_00_15,
    m2.putRq_infoRam_00_14, m3.putRq_infoRam_00_13, m4.putRq_infoRam_00_12,
    m5.putRq_infoRam_00_11, m6.putRq_infoRam_00_10, m7.putRq_infoRam_00_9,
    m8.putRq_infoRam_00_8, m9.putRq_infoRam_00_7, m10.putRq_infoRam_00_6,
    m11.putRq_infoRam_00_5, m12.putRq_infoRam_00_4, m13.putRq_infoRam_00_3,
    m14.putRq_infoRam_00_2, m15.putRq_infoRam_00_1, m16.putRq_infoRam_00_0,
    m17.getRs_dataRam_00, m17.putRq_dataRam_00, m1.getRs_infoRam_00_15,
    m2.getRs_infoRam_00_14, m3.getRs_infoRam_00_13, m4.getRs_infoRam_00_12,
    m5.getRs_infoRam_00_11, m6.getRs_infoRam_00_10, m7.getRs_infoRam_00_9,
    m8.getRs_infoRam_00_8, m9.getRs_infoRam_00_7, m10.getRs_infoRam_00_6,
    m11.getRs_infoRam_00_5, m12.getRs_infoRam_00_4, m13.getRs_infoRam_00_3,
    m14.getRs_infoRam_00_2, m15.getRs_infoRam_00_1, m16.getRs_infoRam_00_0);

    Module64 m64 <- mkModule64 (m27.enq_fifo0002, m38.enq_fifo0012,
    m49.enq_fifo0022, m60.enq_fifo0032, enq_fifo001, enq_fifo000);
    Module65 m65 <- mkModule65 (m19.putRq_infoRam_000_3,
    m20.putRq_infoRam_000_2, m21.putRq_infoRam_000_1,
    m22.putRq_infoRam_000_0, m23.getRs_dataRam_000, m23.putRq_dataRam_000,
    m19.getRs_infoRam_000_3, m20.getRs_infoRam_000_2,
    m21.getRs_infoRam_000_1, m22.getRs_infoRam_000_0);
    Module66 m66 <- mkModule66 (m29.enq_fifo00002, m26.enq_fifo0001,
    m25.enq_fifo0000);
    Module67 m67 <- mkModule67 (m30.putRq_infoRam_001_3,
    m31.putRq_infoRam_001_2, m32.putRq_infoRam_001_1,
    m33.putRq_infoRam_001_0, m34.getRs_dataRam_001, m34.putRq_dataRam_001,
    m30.getRs_infoRam_001_3, m31.getRs_infoRam_001_2,
    m32.getRs_infoRam_001_1, m33.getRs_infoRam_001_0);
    Module68 m68 <- mkModule68 (m40.enq_fifo00102, m37.enq_fifo0011,
    m36.enq_fifo0010);
    Module69 m69 <- mkModule69 (m41.putRq_infoRam_002_3,
    m42.putRq_infoRam_002_2, m43.putRq_infoRam_002_1,
    m44.putRq_infoRam_002_0, m45.getRs_dataRam_002, m45.putRq_dataRam_002,
    m41.getRs_infoRam_002_3, m42.getRs_infoRam_002_2,
    m43.getRs_infoRam_002_1, m44.getRs_infoRam_002_0);
    Module70 m70 <- mkModule70 (m51.enq_fifo00202, m48.enq_fifo0021,
    m47.enq_fifo0020);
    Module71 m71 <- mkModule71 (m52.putRq_infoRam_003_3,
    m53.putRq_infoRam_003_2, m54.putRq_infoRam_003_1,
    m55.putRq_infoRam_003_0, m56.getRs_dataRam_003, m56.putRq_dataRam_003,
    m52.getRs_infoRam_003_3, m53.getRs_infoRam_003_2,
    m54.getRs_infoRam_003_1, m55.getRs_infoRam_003_0);
    Module72 m72 <- mkModule72 (m62.enq_fifo00302, m59.enq_fifo0031,
    m58.enq_fifo0030);
    Module73 m73 <- mkModule73 (m63.cache_00_writeRs,
    m63.cache_00_removeVictim, m63.cache_00_getVictim, m18.transferUpDown00,
    m18.releaseDL00, m18.releaseUL00, m18.upLockGet00, m59.deq_fifo0031,
    m48.deq_fifo0021, m37.deq_fifo0011, m18.addRs00, m18.downLockGet00,
    m26.deq_fifo0001, m64.broadcast_parentChildren00, m18.registerDL00,
    m18.registerUL00, m63.cache_00_hasVictimSlot,
    m64.makeEnq_parentChildren00, m63.cache_00_writeRq, m18.downLockable00,
    m18.upLockable00, m63.cache_00_readRs, m58.deq_fifo0030,
    m47.deq_fifo0020, m36.deq_fifo0010, m25.deq_fifo0000,
    m18.downLockRssFull00, m63.cache_00_readRq, deq_fifo002);
    Module74 m74 <- mkModule74 (m65.cache_000_writeRs,
    m65.cache_000_removeVictim, m65.cache_000_getVictim, m24.releaseUL000,
    m65.cache_000_writeRq, m24.upLockGet000, m24.registerUL000,
    m65.cache_000_hasVictimSlot, m66.makeEnq_parentChildren000,
    m24.downLockable000, m24.upLockable000, m65.cache_000_readRs,
    m28.deq_fifo00000, m24.downLockRssFull000, m65.cache_000_readRq,
    m27.deq_fifo0002);
    Module75 m75 <- mkModule75 (m67.cache_001_writeRs,
    m67.cache_001_removeVictim, m67.cache_001_getVictim, m35.releaseUL001,
    m67.cache_001_writeRq, m35.upLockGet001, m35.registerUL001,
    m67.cache_001_hasVictimSlot, m68.makeEnq_parentChildren001,
    m35.downLockable001, m35.upLockable001, m67.cache_001_readRs,
    m39.deq_fifo00100, m35.downLockRssFull001, m67.cache_001_readRq,
    m38.deq_fifo0012);
    Module76 m76 <- mkModule76 (m69.cache_002_writeRs,
    m69.cache_002_removeVictim, m69.cache_002_getVictim, m46.releaseUL002,
    m69.cache_002_writeRq, m46.upLockGet002, m46.registerUL002,
    m69.cache_002_hasVictimSlot, m70.makeEnq_parentChildren002,
    m46.downLockable002, m46.upLockable002, m69.cache_002_readRs,
    m50.deq_fifo00200, m46.downLockRssFull002, m69.cache_002_readRq,
    m49.deq_fifo0022);
    Module77 m77 <- mkModule77 (m71.cache_003_writeRs,
    m71.cache_003_removeVictim, m71.cache_003_getVictim, m57.releaseUL003,
    m71.cache_003_writeRq, m57.upLockGet003, m57.registerUL003,
    m71.cache_003_hasVictimSlot, m72.makeEnq_parentChildren003,
    m57.downLockable003, m57.upLockable003, m71.cache_003_readRs,
    m61.deq_fifo00300, m57.downLockRssFull003, m71.cache_003_readRq,
    m60.deq_fifo0032);

    //// Initialization logic

    Reg#(Bool) init <- mkReg(False);

    Reg#(Bool) llInitDone <- mkReg(False);
    Reg#(Bit#(10)) llInitIndex <- mkReg(0);

    Reg#(Bool) l1InitDone0 <- mkReg(False);
    Reg#(Bit#(8)) l1InitIndex0 <- mkReg(0);
    Reg#(Bool) l1InitDone1 <- mkReg(False);
    Reg#(Bit#(8)) l1InitIndex1 <- mkReg(0);
    Reg#(Bool) l1InitDone2 <- mkReg(False);
    Reg#(Bit#(8)) l1InitIndex2 <- mkReg(0);
    Reg#(Bool) l1InitDone3 <- mkReg(False);
    Reg#(Bit#(8)) l1InitIndex3 <- mkReg(0);

    function Struct22 llDefaultLine (Bit#(49) tagValue);
      return Struct22 { write: True,
                       addr: llInitIndex,
                       datain: Struct19 { tag: tagValue,
                                         value: Struct4 { mesi_owned: False,
                                                         mesi_status: 3'h1,
                                                         mesi_dir_st: 3'h1,
                                                         mesi_dir_sharers: 4'h0 }}};
    endfunction

    rule ll_info_do_init (!llInitDone);
        m1.putRq_infoRam_00_15 (llDefaultLine(15));
        m2.putRq_infoRam_00_14 (llDefaultLine(14));
        m3.putRq_infoRam_00_13 (llDefaultLine(13));
        m4.putRq_infoRam_00_12 (llDefaultLine(12));
        m5.putRq_infoRam_00_11 (llDefaultLine(11));
        m6.putRq_infoRam_00_10 (llDefaultLine(10));
        m7.putRq_infoRam_00_9 (llDefaultLine(9));
        m8.putRq_infoRam_00_8 (llDefaultLine(8));
        m9.putRq_infoRam_00_7 (llDefaultLine(7));
        m10.putRq_infoRam_00_6 (llDefaultLine(6));
        m11.putRq_infoRam_00_5 (llDefaultLine(5));
        m12.putRq_infoRam_00_4 (llDefaultLine(4));
        m13.putRq_infoRam_00_3 (llDefaultLine(3));
        m14.putRq_infoRam_00_2 (llDefaultLine(2));
        m15.putRq_infoRam_00_1 (llDefaultLine(1));
        m16.putRq_infoRam_00_0 (llDefaultLine(0));

        llInitIndex <= llInitIndex + 1;
        if (llInitIndex == maxBound) begin
            llInitDone <= True;
        end
    endrule

    function Struct29 l1DefaultLine (Bit#(51) tagValue, Bit#(8) index);
      return Struct29 { write: True,
                       addr: index,
                       datain: Struct26 { tag: tagValue,
                                         value: Struct4 { mesi_owned: False,
                                                         mesi_status: 3'h1,
                                                         mesi_dir_st: 3'h1,
                                                         mesi_dir_sharers: 4'h0 }}};
    endfunction

    rule l1_info_do_init_0 (!l1InitDone0);
        m19.putRq_infoRam_000_3 (l1DefaultLine(3, l1InitIndex0));
        m20.putRq_infoRam_000_2 (l1DefaultLine(2, l1InitIndex0));
        m21.putRq_infoRam_000_1 (l1DefaultLine(1, l1InitIndex0));
        m22.putRq_infoRam_000_0 (l1DefaultLine(0, l1InitIndex0));
        l1InitIndex0 <= l1InitIndex0 + 1;
        if (l1InitIndex0 == maxBound) begin
            l1InitDone0 <= True;
        end
    endrule

    rule l1_info_do_init_1 (!l1InitDone1);
        m30.putRq_infoRam_001_3 (l1DefaultLine(3, l1InitIndex1));
        m31.putRq_infoRam_001_2 (l1DefaultLine(2, l1InitIndex1));
        m32.putRq_infoRam_001_1 (l1DefaultLine(1, l1InitIndex1));
        m33.putRq_infoRam_001_0 (l1DefaultLine(0, l1InitIndex1));
        l1InitIndex1 <= l1InitIndex1 + 1;
        if (l1InitIndex1 == maxBound) begin
            l1InitDone1 <= True;
        end
    endrule

    rule l1_info_do_init_2 (!l1InitDone2);
        m41.putRq_infoRam_002_3 (l1DefaultLine(3, l1InitIndex2));
        m42.putRq_infoRam_002_2 (l1DefaultLine(2, l1InitIndex2));
        m43.putRq_infoRam_002_1 (l1DefaultLine(1, l1InitIndex2));
        m44.putRq_infoRam_002_0 (l1DefaultLine(0, l1InitIndex2));
        l1InitIndex2 <= l1InitIndex1 + 1;
        if (l1InitIndex2 == maxBound) begin
            l1InitDone2 <= True;
        end
    endrule

    rule l1_info_do_init_3 (!l1InitDone3);
        m52.putRq_infoRam_003_3 (l1DefaultLine(3, l1InitIndex3));
        m53.putRq_infoRam_003_2 (l1DefaultLine(2, l1InitIndex3));
        m54.putRq_infoRam_003_1 (l1DefaultLine(1, l1InitIndex3));
        m55.putRq_infoRam_003_0 (l1DefaultLine(0, l1InitIndex3));
        l1InitIndex3 <= l1InitIndex1 + 1;
        if (l1InitIndex3 == maxBound) begin
            l1InitDone3 <= True;
        end
    endrule

    rule init_done (!init && llInitDone &&
                    l1InitDone0 && l1InitDone1 && l1InitDone2 && l1InitDone3);
        init <= True;
    endrule

    function MemRqRs getMemRqRs (function Action enq_rq (Struct2 _),
                                 function ActionValue#(Struct2) deq_rs ());
        return interface MemRqRs;
                   method mem_enq_rq = enq_rq;
                   method mem_deq_rs = deq_rs;
               endinterface;
    endfunction

    Vector#(L1Num, MemRqRs) _l1Ifc = newVector();
    _l1Ifc[0] = getMemRqRs(m28.enq_fifo00000, m29.deq_fifo00002);
    _l1Ifc[1] = getMemRqRs(m39.enq_fifo00100, m40.deq_fifo00102);
    _l1Ifc[2] = getMemRqRs(m50.enq_fifo00200, m51.deq_fifo00202);
    _l1Ifc[3] = getMemRqRs(m61.enq_fifo00300, m62.deq_fifo00302);
    interface l1Ifc = _l1Ifc;

    interface DMA llDma;
        method dma_putRq = m17.putRq_dataRam_00;
        method dma_getRs = m17.getRs_dataRam_00;
    endinterface

    method Bool isInit ();
        return init;
    endmethod

endmodule
